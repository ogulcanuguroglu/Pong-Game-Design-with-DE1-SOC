library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity main is
  port(
      CLOCK_50, RST: in STD_LOGIC;
		SW2 : in STD_LOGIC;
		p1_up, p1_down : in std_logic;
		p2_up, p2_down : in std_logic;
      VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_N, VGA_SYNC_N: out STD_LOGIC;
      VGA_R, VGA_G, VGA_B: out STD_LOGIC_VECTOR(7 downto 0) --8 pins for RGB
      );
end entity main;

architecture rtl of main is

    constant HD  : integer   := 640; --  640   Horizontal Display (640)
    constant HFP : integer   := 16;  --   16   Right border (front porch)
    constant HSP : integer   := 96;  --   96   Sync pulse (Retrace)
    constant HBP : integer   := 48;  --   48   Left boarder (back porch)

    constant VD  : integer   := 480; --  480   Vertical Display (480)
    constant VFP : integer   := 10;  --   10   Right border (front porch)
    constant VSP : integer   := 2;   --    2   Sync pulse (Retrace)
    constant VBP : integer   := 33;  --   33   Left boarder (back porch)
	 
	 constant TOT_H : integer := 800;

	 constant TOT_V : integer := 800;	
    
	 signal clk25 : std_logic := '0';

    signal hPos  : integer   := 0;
    signal vPos  : integer   := 0;

    signal hs    : std_logic := '0'; -- register to account for pixel data delay
    signal vs    : std_logic := '0'; -- register to account for pixel data delay
    signal de    : std_logic := '0';

	 signal ball_x1: integer range 1 to TOT_H := 313;
	 signal ball_x2: integer range 1 to TOT_H := 327;
	 signal ball_y1: integer range 1 to TOT_H := 233;
	 signal ball_y2: integer range 1 to TOT_H := 247;
	 signal ball_move_h: integer range -200 to 200 := 1;
	 signal ball_move_v: integer range -200 to 200 := 1;
	 
	 signal p1_x1: integer range 1 to TOT_H := 20;
	 signal p1_x2: integer range 1 to TOT_H := 32;
	 signal p1_y1: integer range 1 to TOT_H := 195;
	 signal p1_y2: integer range 1 to TOT_H := 285;
	 
	 
	 signal p2_x1: integer range 1 to TOT_H := 608;
	 signal p2_x2: integer range 1 to TOT_H := 620;
	 signal p2_y1: integer range 1 to TOT_V := 195;
	 signal p2_y2: integer range 1 to TOT_V := 285;

	 
	 signal delayCounter1, delayCounter2, delayCounter3 : integer range 0 to 100000;
	 
	 signal newGame : std_logic;
	 signal gameLabelVisible, logoVisible : std_logic;
	 signal label_0p1_visible: std_logic;
	 signal label_1p1_visible: std_logic;
	 signal label_2p1_visible : std_logic;	 
	 signal label_3p1_visible: std_logic;
	 signal label_0p2_visible: std_logic;
	 signal label_1p2_visible: std_logic;
	 signal label_2p2_visible : std_logic;	 
	 signal label_3p2_visible: std_logic;
	 signal P1_Won_Label_visible: std_logic;	 
	 signal P2_Won_Label_visible: std_logic;	 
	 signal StartGameLabelVisible: std_logic;
	 
	 type BITMAP1 is array (0 to 173) of std_logic_vector(0 to 399);
	 type BITMAP2 is array (0 to 46) of std_logic_vector(0 to 399);
	 type BITMAP3 is array (0 to 164) of std_logic_vector(0 to 199);
	 type BITMAP4 is array (0 to 63) of std_logic_vector(0 to 399);
	 type BITMAP5 is array (0 to 63) of std_logic_vector(0 to 399); 
	 type BITMAP6 is array (0 to 103) of std_logic_vector(0 to 83);
	 type BITMAP9 is array (0 to 48) of std_logic_vector(0 to 399);
	 
	 type BITMAP7 is array (0 to 13) of std_logic_vector(0 to 78);
	 signal p1_label: BITMAP7;
	 signal p1_label_visible : std_logic;
	 signal p2_label: BITMAP7;
	 signal p2_label_visible : std_logic;
	 
		
	 signal label_0: BITMAP6;
	 signal label_1: BITMAP6;
	 signal label_2: BITMAP6;
	 signal label_3: BITMAP6;
	 signal P1_Won_Label: BITMAP1;
	 signal P2_Won_Label: BITMAP1;
	 signal StartGameLabel: BITMAP9;
	 
	 signal logo: BITMAP3;
	 signal gameLabel: BITMAP4;
	 
	 type g_State is (MENU, INITIAL, GAME, P1_WIN, P2_WIN);
	 signal current_state, next_state: g_State := MENU;
	 signal p1_w, p2_w : std_logic;
	 
	 signal score_p1 : integer := 0;
	 signal score_p2 : integer := 0;
	 
	 signal delay_label : integer := 0;	 
	 signal goal_flag : std_logic := '0';
	 signal label_delay_on : std_logic;
	 
begin
p1_label <=(
"1111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1100000000111000011111111111111111111111111111111111111111111111111111000111111",
"1100111100011110011111111111111111111111111111111111111111111111111100000111111",
"1100111100011110011111100000011100111110011110000001110001000011111110000111111",
"1100111100011110011111100000001100011110001100000001110001000011111111000111111",
"1100111100011110011111111111000100011110001000111100010000111111111111000111111",
"1100000000111110011111100000000100011110001000000000010001111111111111000111111",
"1100000000111110011111000000000100000000001000000000110001111111111111000111111",
"1100111111111110001110001111000110000000001000111111110001111111111111000111111",
"1100111111110000000011100000000111111110001100000001110001111111111000000001111",
"1111111111111111111111111111111110000000111111111111111111111111111111111111111",
"1111111111111111111111111111111111000000111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111"
);

p2_label <=(
"1111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1100000000111000011111111111111111111111111111111111111111111111111111000111111",
"1100111100011110011111111111111111111111111111111111111111111111111110000001111",
"1100111100011110011111100000011100111110011110000001110001000011111110011001111",
"1100111100011110011111100000001100011110001100000001110001000011111111111001111",
"1100111100011110011111111111000100011110001000111100010000111111111111110011111",
"1100000000111110011111100000000100011110001000000000010001111111111111100011111",
"1100000000111110011111000000000100000000001000000000110001111111111111000111111",
"1100111111111110001110001111000110000000001000111111110001111111111110001111111",
"1100111111110000000011100000000111111110001100000001110001111111111110000001111",
"1111111111111111111111111111111110000000111111111111111111111111111110000001111",
"1111111111111111111111111111111111000000111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111"
);

gameLabel <= ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111000000000000000000000011111111111111111111111111111111000000011111111111111111111111111111111110000000000011111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111100000000001111111111111111111111111111111000000000011111111110000000000111111111111111111111111111111100000000000111111111111111111111111",
                  "1111111011111111111111111100000111111111111111111111111110000000000000011111111111111111111111111111000001111100000111111111111111111111111111100000111110000011111111111111111111111111111111111111111111111111111111111100000111100000011111111111111111111111111100000011111000001111111111111111111111111100000111110000111111000001111100000111111111111111111111111100000011111000001111111111111111111111",
                  "1111111011111111111111111111110001111111111111111111111000011111111110000111111111111111111111111100001111111111110001111111111111111111111110001111111111110000111111111111111111111111111111111111111111111111111111110001111111111110001111111111111111111111110000111111111111000111111111111111111111110001111111111110001100011111111111100011111111111111111111111000111111111111000011111111111111111111",
                  "1111111011000000000000000000011100111111111111111111110001111000000011110001111111111111111111111000111000000000011100111111111111111111111100011100000000111100011111111111111111111111111111111111111111111111111111000111100000000111100111111111111111111111100011100000000001110001111111111111111111100111000000000011100001110000000000111001111111111111111111100011100000000001110001111111111111111111",
                  "1111111011011111111111111110000110011111111111111111100111100000000000011000111111111111111111110011100001111110000110001111111111111111111001110000011100000110001111111111111111111111111111111111111111111111111110001110000111100001110001111111111111111111000110000111111000011100111111111111111111001100001111110000110011000011111100001100111111111111111111000110000111111000011100111111111111111111",
                  "1111111011011111111111111111100011001111111111111111001110011111111111001110011111111111111111100110001111111111100011000111111111111111110011000111111111100011000111111111111111111111111111111111111111111111111100011000111111111100011000111111111111111110011100111111111111001110011111111111111110011000111111111100011110001111111111000110011111111111111110011100011111111111001110011111111111111111",
                   "1111111011011000000000000000111001100111111111111110011100111000000011100011001111111111111111001100111100000000111001100111111111111111100110011110000000111001100011111111111111111111111111111111111111111111111000110011110000001111001100111111111111111100111001110000000011100011001111111111111110110001110000000111001100011000000001110011001111111111111100111001110000000011100011001111111111111111",
                  "1111111011011001111111111100001100110011111111111100111011100000000000111001100111111111111110011001110000111100001100110011111111111111001100111000000000001100110001111111111111111111111111111111111111111111111001100110000000000001100110011111111111111100110011000011110000110011000111111111111100100011000011100011100001110001111000111001100111111111111100110011000011110000111001100111111111111111",
                  "1111111011011011111111111111000110011001111111111100110010000111111110001100110011111111111110010011000111111111000110011001111111111110011001100011111111100110011000111111111111111111111111111111111111111111110011001100011111111000110011001111111111111001100110011111111110011001100011111111111101100110001111111001110001100111111110011100100011111111111001100110011111111110011101110011111111111111",
                  "1111111011011011000000000001110011001000111111111001100100011100000111000110110001111111111100110010001100000001110011001000111111111110010011000110000001110011001100011111111111111111111111111111111111111111110110011001110000001110011001000111111111110011001100110000000111001100110001111111111001001100110000001100110011001100000011001100110001111111111011001100111000000011001100110001111111111111",
                  "1111111011011011000000000000011001001100011111111001001100110000000001100010011000111111111100100110010000000000011001001100011111111100110010001100000000011001100100001111111111111111111111111111111111111111100110110011000000000011001001100011111111110010011001100000000001100110010000111111111001001100100000000110011010011000000001100110110000111111110011011001100000000001100110011000111111111111",
                  "1111111011011011000000000000001001100100001111110011001001100000000000010011001000011111111001101100100000000000001001100100001111111100100110010000000000001100100110000111111111111111111111111111111111111111101100100110000000000001101100100001111111110110010011000000000000110010011000011111111011001001100000000010011110010000000000100110010000011111110010011011000000000000110011011000011111111111",
                  "1111111011011011000000000000000100100100000111110010011001000000000000011001001000001111111001001101100000000000001100100110000111111101100100110000000000000110110010000111111111111111111111111111111111111111001101100100000000000000100100110000111111100110110010000000000000010011011000011111111011011001000000000011001110110000000000110010010000011111110110010010000000000000011011001000001111111111",
                  "1111111011011011000000000000000100110110000111110010010011000000000000001001101100001111111001001001000000000000000100110110000011111101101100100000000000000110010010000011111111111111111111111111111111111111001001101100000000000000110110010000011111100100110110000000000000011011001000001111110011011011000000000001001100100000000000010010010000001111100110110110000000000000011001001000001111111111",
                  "1111111011011011000000000000000110110110000011110110010010000000000000001101101100000111111011001001000000000000000110110010000011111001101100100000000000000010010010000001111111111111111111111111111111111111001001001100000000000000110010010000011111100100100100000000000000001001001000001111110011011011000000000001001100100000000000010010010000001111100100100110000000000000001001001100000111111111",
                  "1111111011011011000000000000000010110010000001110110110010000000000000001101100100000111111011011001000000000000000110110010000001111001001101100000000000000011011011000001111111111111111111111111111111111111001001001000000000000000010010010000001111100100100100000000000000001001001000000111110011011011000000000001101101100000000000010010011000000111100100100100000000000000001001101100000111111111",
                  "1111111011011011000000011111110010110010000001110110110010000000000111101101100100000011111011011001000000000111110110110010000001111001001101100000000001110010011011000000111111111111111111111111111111111111001001001000000000011110010010010000001111100100100100000000001111001001001000000111110011011011000000001101101101100000000010010010011000000111100100100100000000001111001001101100000011111111",
                  "1111111011011011000000011111110010110010000001110110110010000000011111101101100100000011111011011001000000001111110110110010000001111001001101100000000111110000000000000000111111111111111111111111111111111111001001001000000000111110000000000000000111100100100100000000011111001001001000000011110011011011000000011101101101100000000110010010011000000111100100100100000000011111000000000000000011111111",
                  "1111111011011011000000011111100110110110000001110110110010000000011111101101100100000011111011011001000000001111110110110010000000111001001101100000001111111000000000000000111111111111111111111111111111111111001001001000000001111110000000000000000111100100100100000000111111001001001000000011110011011011000000011101101101100000001110010010011000000111100100100100000000111111100000000000000011111111",
                  "1111111011011011000000011111100100110110000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111100000000000000111111111111111111111111111111111111001001001000000001111111100000000000000111100100100100000001111111001001001000000011110011011011000000011101101101100000001110010010011000000111100100100100000000111111110000000000000011111111",
                  "1111111011011011000000011111100100100110000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111110000000000000111111111111111111111111111111111111001001001000000011111111110000000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111111000000000000011111111",
                  "1111111011011011000000011111001001100100000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111111111000000000000111111111111111111111111111111111111001001001000000011111111111000000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111111100000000000001111111",
                  "1111111011011011000000011100011001101100000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111100000000000111111111111111111111111111111111111001001001000000011111111111000000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111111110000000000001111111",
                  "1111111011011011000000000001110011001000000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000000000000000111111111111111111111111111111111111001001001000000000000000000000000000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000011111000000000011111111",
                  "1111111011011011111111111111000110011000000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111111111000111111111111111111111111111111111111111001001001000000001111111111111110001111111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111111001111111111111111111111",
                  "1111111011011001111111111100001100110000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111111111000011111111111111111111111111111111111111001001001000000001111111111111110000111111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111111000111111111111111111111",
                  "1111111011011000000000000000111001100000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000000011000001111111111111111111111111111111111111001001001000000000000000000000010000011111100100100000000000000000000001001000000011110011011011000000111101101101100000001110010010011000000111100100100000000000000000000011111111111111111111",
                  "1111111011011111111111111111100011100000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000000011000000111111111111111111111111111111111111001001001000000000000000000000010000001111100100111111111111111111111111001000000011110011011011000000111101101101100000001110010010011000000111100100111111111111111110000000111111111111111111",
                  "1111111011011111111111111110000110000000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111111011000000111111111111111111111111111111111111001001001000000001111111111110010000000111100100111111111111111111111111001000000011110011011011000000111101101101100000001110010010011000000111100100111111111111111111000000111111111111111111",
                  "1111111011011000000000000000011100000000000011110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000011011000000111111111111111111111111111111111111001001001000000000000000000010010000000111100100100000000000000000000001001000000011110011011011000000111101101101100000001110010010011000000111100100100000000000000000000000111111111111111111",
                  "1111111011011001111111111111110000000000000011110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000011011000000111111111111111111111111111111111111001001001000000000000000000010010000000111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111110000000111111111111111111",
                  "1111111011011011111111111110000000000000000111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111011011000000111111111111111111111111111111111111001001001000000001111111110010010000000111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111111000000111111111111111111",
                  "1111111011011011000000000000000000000000001111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000011011011000000111111111111111111111111111111111111001001001000000000000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000000011111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000011011011000000111111111111111111111111111111111111001001001000000000000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000000111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000011011011000000111111111111111111111111111111111111001001001000000010000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000001111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011000000011011011000000111111111111111111111111111111111111001001001000000011000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011100000011011011000000111111111111111111111111111111111111001001001000000011100000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000011111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011110000011011011000000111111111111111111111111111111111111001001001000000011110000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000011111111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111000011011011000000111111111111111111111111111111111111001001001000000011111000010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000000000111111111111",
                  "1111111011011011000000011111111111111111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111110011011011000000111111111111111111111111111111111111001001001000000011111110010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111001000000100011111111111",
                  "1111111011011011000000011111111111111111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111110011011011000000111111111111111111111111111111111111001001001000000011111110010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111001101101100001111111111",
                  "1111111011011011000000011111111111111111111111110110010010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111110010011011000000111111111111111111111111111111111111001001001000000011111110010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100110000001111111011001101100000111111111",
                  "1111111011011011000000011111111111111111111111110010010011000000111111001001101100000001111011011001000000011111110110110010000000111001101100100000011111110010010010000000111111111111111111111111111111111111001001101100000011111110110010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100110110000001111110011001001100000011111111",
                  "1111111011011011000000011111111111111111111111110010011011000000111111001001001100000001111011011001000000011111110110110010000000111101100100100000011111110110010010000000111111111111111111111111111111111111001101100100000011111100110110010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100110110010000001111110011001001000000011111111",
                  "1111111011011011000000011111111111111111111111110011001001100000111110011011001000000001111011011001000000011111110110110010000000111100100110110000011111100100110010000000111111111111111111111111111111111111101100100110000011111000100110110000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111110110010011000001111100110011011000000001111111",
                  "1111111011011011000000011111111111111111111111111011001001110000111000010011011000000001111011011001000000011111110110110010000000111100110110011000011110001100100110000000111111111111111111111111111111111111100100110010000011110001000100100000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111110010011001100001110001110010011000000001111111",
                  "1111111011011011000000011111111111111111111111111001100100111000000001100110011000000001111011011001000000011111110110110010000000111110010011001100000000011001100100000000111111111111111111111111111111111111100110011001100000000010001101100000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111110011001100110000000011100110110000000001111111",
                  "1111111011011011000000011111111111111111111111111001100110011110001111001100110000000001111011011001000000011111110110110010000000111110011001100111100011110011001100000000111111111111111111111111111111111111110010001000111100011100011001000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111001100110001111111110001100110000000011111111",
                  "1111111011011011000000011111111111111111111111111100110011000111111100011100100000000001111011011001000000011111110110110010000000111111001100110001111111000110011000000000111111111111111111111111111111111111110011001110001111110000110011000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111100100011000001111000011001100000000011111111",
                  "1111111011011011000000011111111111111111111111111110011001100000000000111001100000000011111011011001000000011111110110110010000000111111000110011100000000001100010000000000111111111111111111111111111111111111111001100011000000000001100110000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111100110001110000000001110011000000000011111111",
                  "1111111011011011000000011111111111111111111111111110001100011100000111100011000000000011111011011001000000011111110110110010000000111111100011001111000001111000100000000000111111111111111111111111111111111111111100110001111000001110001100000000001111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111110011100111111111111000110000000000011111111",
                  "1111111011011011000000011111111111111111111111111111000110001111111110001110000000000011111011011001000000011111110110110010000000111111110001100011111111100011000000000001111111111111111111111111111111111111111110011100011111111000011000000000001111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111000110000111111100011100000000000111111111",
                  "1111111011011011000000011111111111111111111111111111100011100000000000011100000000000111111011011001000000011111110110110010000000111111111000111000000000000110000000000001111111111111111111111111111111111111111111000110000000000001110000000000001111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111100011100000000001111000000000000111111111",
                  "1111111011011011000000011111111111111111111111111111110001111000000011110000000000000111111011011001000000011111110110110010000000111111111100011111000001111100000000000011111111111111111111111111111111111111111111100011110000001111000000000000011111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111110000111111111111100000000000001111111111",
                  "1111111011011011000000011111111111111111111111111111111100001111111111000000000000001111111011011001000000011111110110110010000000111111111110000011111111100000000000000011111111111111111111111111111111111111111111110000111111111100000000000000111111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111111000000111111100000000000000001111111111",
                  "1111111000000000000000011111111111111111111111111111111110000000000000000000000000011111111000000000000000011111110000000000000000111111111111000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000111111100000000000000001111111000000000000000011110000000000000000111100000000000000001110000000000000000111111111111100000000000000000000000000011111111111",
                  "1111111000000000000000011111111111111111111111111111111111000000000000000000000000011111111000000000000000011111110000000000000000111111111111100000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000001111111100000000000000001111111000000000000000011111000000000000000111100000000000000001110000000000000000111111111111110000000000000000000000000111111111111",
                  "1111111100000000000000011111111111111111111111111111111111100000000000000000000000111111111100000000000000011111111000000000000000111111111111110000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000011111111110000000000000001111111110000000000000011111100000000000000111110000000000000001111100000000000000111111111111111100000000000000000000001111111111111",
                  "1111111110000000000000011111111111111111111111111111111111110000000000000000000011111111111110000000000000011111111100000000000000111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111000000000000000000000111111111111000000000000001111111111000000000000011111110000000000000111111000000000000001111110000000000000111111111111111110000000000000000000011111111111111",
                  "1111111111000000000000011111111111111111111111111111111111111000000000000000000111111111111111000000000000011111111110000000000000111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000011111111111111100000000000001111111111100000000000011111111000000000000111111100000000000001111111000000000000111111111111111111000000000000000001111111111111111",
                  "1111111111100000000000011111111111111111111111111111111111111110000000000000011111111111111111100000000000011111111111000000000000111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000001111111111110000000000011111111100000000000111111110000000000001111111100000000000111111111111111111110000000000000111111111111111111",
                  "1111111111110000000000111111111111111111111111111111111111111111100000000011111111111111111111110000000000111111111111100000000000111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111100000000001111111111111000000000011111111110000000000111111111000000000011111111110000000000111111111111111111111111000001111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
    --The process involves the next state logic for the variables
logo <= (	 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111100000000001100000000000001111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111100000000011000000000000111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111110000000011000000000001111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111000000011100000000001111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000001110000000001111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111110000001110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111000000111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111100000011110000000001111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111000001111000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111100000011100000000011111111111111111111111111111111111111111111111111111111111111111111111111000001000010000100000001111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111000001111000000001111111111111111111111111111111111111111111111111111111111111111111111111000010000000010001111111000011111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111100000011100000000011111111111111111111111111111111111111111111111111111111111111111111111100000010000100111111110011000000111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111000001111000000001111111111111111111111111111111111111111111111111111111111111111111111111000000011001111111000100001000100001111111111111111111111111111",
             "11111111111111111111111111111111111111111111110000011110000000011111111111111111111111111111111111111111111111111111111111111111111111100000110111101110001000100001100111000111111111111111111111111111",
             "11111111111111111111111111111111111111111111100001111000000001111111111111111111111111111111111111111111111111111111111111111111111111000111110011000100001000110011111111000011111111111111111111111111",
             "11111111111111111111111111111111111111111110000011110000000011111111111111111111111111111111111111111111111111111111111111111111111100011000100001000000001101111111100010001000111111111111111111111111",
             "11111111111111111111111111111111111111111100000111100000000111111111111111111111111111111111111111111111111111111111111111111111111000001000100001000111111110110001100010001100011111111111111111111111",
             "11111111111111111111111111111111111111111000001111000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000110011111111001100010000100011111110001111111111111111111111",
             "11111111111111111111111111111111111111110000011110000000111111111111111111111111111111111111110000000001111111111111111111111111100000001000111111100010000100011001111111111110000111111111111111111111",
             "11111111111111111111111111111111111111100001111100000001111111111111111111111111111111111111000000000000111111111111111111111111000110011110110001000010000100011111111111000110000111111111111111111111",
             "11111111111111111111111111111111111111000011111000000011111111111111111111111111111111111111000000000000111111111111111111111110001111001100010000100011001111111100110001000110010011111111111111111111",
             "11111111111111111111111111111111111110000111110000000111111111111111111111111111101111111111000000000000011111111111111111111100100010000000010000110111111110011000110001100111111001111111111111111111",
             "11111111111111111111111111111111111100001111100000001111111111111111111111111110000111111111000001100000011111111111111111111000000010000100011111111011000100001000110011111111111101111111111111111111",
             "11111111111111111111111111111111111000011111000000011111111111111111111111111000000111111111000001100000011111111111111111110000000010001111111100100001000110001101111111110111001100111111111111111111",
             "11111111111111111111111111111111111000111110000000011111111111111111111111111100000011111111000001111111111111111111111111100000100011111110001000000001000111111111111001100011001110011111111111111111",
             "11111111111111111111111111111111110000111100000000111111111111111111111111111100000011111111000001111111111111111111111111001001111011000100001000010001111111111100010001100011111110011111111111111111",
             "11111111111111111111111111111111100001111000000001111111111111111111111000011110000001111111000001111111111111111111111110011100100001000000001100111111110110001100011001111111111111001111111111111111",
             "11111111111111111111111111111111000011110000000011111111111111111111100000001110000001111111000001000000011111111111111110001000100001000110011111111001100010000100011111111111101110001111111111111111",
             "11111111111111111111111111111110000111110000000111111111111111111111110000000111000000111111000001100000011111111111111100001000010001101111111100010000100011001111111111110011100111000111111111111111",
             "11111111111111111111111111111110001111100000001111111111111111111111110000000001000000111111000001100000011111111111111000001000111111100010000100010000110111111111011000110011101111100111111111111111",
             "11111111111111111111111111111100001111000000001111111111111111111111111000000000100000011111000001110000011111111111111000001111111001100010000100011111111111100110001000111011111111110111111111111111",
             "11111111111111111111111111111000011110000000011111111111111111111111111000000000000000011111000001110000011111111111110011111100010000100010001111111111110001000110001111111111111111000011111111111111",
             "11111111111111111111111111110000111110000000111111111111111111111111111100000000000000001111000000110000011111111111110010000000010000100011111110011000110001000111111111111111100111000011111111111111",
             "11111111111111111111111111110001111100000000111111111111111111011111111100000000000000001111000000110000011111111111100010000100011001111111000110001000110011111111111110111001110111110011111111111111",
             "11111111111111111111111111100001111000000001111111111111111110001111111110000000000000000111000000110000011111111111100000000110111101110001000010001100111111111111001100011001111111111011111111111111",
             "11111111111111111111111111100011111000000001111111111111111100000111111110000000000000000111000000000000001111111111000011111110011000100001000110011111111001100011001100111111111111111011111111111111",
             "11111111111111111111111111000111110000000011111111111111111000000011111111000000000000000011100000000000001111111111011111100110001000010001101111111100011000100011001111111111111111100001111111111111",
             "11111111111111111111111110000111110000000111111111111111111100000001111111000000110000000011100000000000001111111111010001000000001000111111111111001100011000110111111111111100110011101001111111111111",
             "11111111111111111111111110001111100000000111111111111111111110000000111111100000011000000001111000001111111111111110000001000010001111111001100010000100011111111111101110011100111111111001111111111111",
             "11111111111111111111111100001111100000001111111111111111111111000000011111100000011110000001111111111111111111111110000001100111111100010000100011001111111111111011100110001111111111111001111111111111",
             "11111111111111111111111100011111000000001111111111111111111111100000001111110000001111000111111111111111111111111110010011111111001100010000100011111111111100110001100111111111111111110001111111111111",
             "11111111111111111111111000011111000000011111111111111111111111110000000111110000001111111111111111111111111111111110111001100010000100011001111111101110001000110011111111111111111001110001111111111111",
             "11111111111111111111111000111110000000011111111111111111111111111000000011111000000111111111111111111111111111111110010000100010000110111111110011000110001100111111111111001110011001111001111111111111",
             "11111111111111111111110000111110000000011111111111111111111111111100000001111000000111111111111111111111111111111110010000100011111111111100110001000111011111111111110011001110111111111001111111111111",
             "11111111111111111111110001111100000000111111111111111111111111111110000000111100001111111111111111111111111111111110011001111111100110001000010001101111111110111001100011101111111111111011111111111111",
             "11111111111111111111100001111100000000111111111111111000011111111111000000011100111111111111111111111111111111111110011111110011000110001000111111111111001100011001111111111111111111111011111111111111",
             "11111111111111111111100011111000000001111111111111110000000111111111100000001111111111111111111111111111111111111110011100110001000110001111111111100011000100011111111111111111011100110011111111111111",
             "11111111111111111111100011111000000001111111111111100000000001111111110000000111111111111111111111111111111111111110001000010001100111111110111000100011001111111111111111100111011111110011111111111111",
             "11111111111111111111000111111000000001111111111111100000000000011111111000000111111111111111111111111111111111111110001000111011111111001100011000110011111111111100110011100111111111110111111111111111",
             "11111111111111111111000111110000000011111111111111000000000000001111111100001111111111111111111111111111111111111111001111111111100011000100011001111111111110011100111011111111111111100111111111111111",
             "11111111111111111110000111110000000011111111111111000011000000000111111110011111111111111111111111000000111111111111001111111000100011000110111111111111100110001100111111111111111110100111111111111111",
             "11111111111111111110001111100000000011111111111110000011110000000111111111111111111111111111111111001110001111111111000100010000100011111111111100110001100111011111111111111111101111101111111111111111",
             "11111111111111111110001111100000000111111111111110000011111100000111111111111111111111111111111110011111100111111111100000011001111111111110001000110001111111111111111101110011111111001111111111111111",
             "11111111111111111100001111100000000111111111111100000000111100001111111111111111111111111111111100111111110011111111100000011111111111100110001100111111111111111110011001111111111111011111111111111111",
             "11111111111111111100011111100000000111111111111100000000001000001111111111111111111111111111111001111111111001111111100100111100110001000110001111111111110111001110011111111111111110011111111111111111",
             "11111111111111111100011111000000000111111111111100000000000000011111111111111111111111111111110011111111111100111111100110001000110001100111111111111001100011001111111111111111111100111111111111111111",
             "11111111111111111000011111000000001111111111111111000000000000011111111111111111111111111111100011111111100110011111100111001100111011111111111110011001110011111111111111111011000000000111111111111111",
             "11111111111111111000111111000000001111111111111111110000000000001111111111111111111111111111100111111111000010011111100111100111111111110111000100011001111111111111111100111000001111000001111111111111",
             "11111111111111111000111111000000001111111111111111111100000000000011111111111111111111111111001111111110000011011111100111110011111001100011001110111111111111100111011111111000111000110000111111111111",
             "11111111111111111000111110000000001111111111111111111111000000000000111111111111111111111110011111111100000001001111100111111000011000110011111111111111111011100111111111110011111100000100011111111111",
             "11111111111111110000111110000000001111111111111111111111110000000000111111111111111111111100111111111000000001001111100111111100011001111111111111011100111011111111111111100111111100000000001111111111",
             "11111111111111110001111110000000001111111111111111111111111100000000111111111111111111111001111111110000000011001111100111111110011111111111100110001100111111111111111111001101111000000000001111111111",
             "11111111111111110001111110000000011111111111111111111111111111000001111111111111111111110011111111100000000110011111101111011111001111110001100111011111111111111111101110001001100000000000000111111111",
             "11111111111111110001111110000000011111111111111111111111111111110001111111111111111111100111111111000000001100111111101110111111100100110001100111111111111111110011101111011000000000000000000111111111",
             "11111111111111110001111100000000011111111111111111111111111111111111111111111111111111000111111110000000111001111111001101101111110000111111111111111110111001110111111110010001110000000000000111111111",
             "11111111111111110001111100000000011111111111111111111111111111111111111111111111111110001111111100000001100011111111000011011111111001111111111111001110011111111111111110010001000000000000000011111111",
             "11111111111111100011111100000000011111111111111111111111111111111111111111111111111100011111111000000011000111111110000111011111111100111111110011001111111111111111111110010000000000000000000011111111",
             "11111111111111100011111100000000011111111111111111111111111111111111111111111111111000111111110000000110011111111110001111011111111110011001110011111111111111111111111110010000000000000000000011111111",
             "11111111111111100010000000000000011111111111111111111111111111111111111111111111110001111111100000001100111111111100011001011111111111001001111111111111111110111011111110010000000000000000000111111111",
             "11111111111111100000000000000000011111111111111111111111111111111111111111111111100111111111000000011001111111111000110001001111110111100111111111111111011110111111111100010000000000000000000111111111",
             "11111111111111100000000000000000011111111111111111111111111111111111111111111111000111111110000001110011111111110001100001100011001111110011111011100111011111111111111000000000000000000000000111111111",
             "11111111111111100001111111110000011111111111111111111111111111111111111111111110011111111100000011000111111111100011000000111000110111111000111001111111111111111111110011001000000000000000000111111111",
             "11111111111111100111111111111100011111111111111111000000001111111111111111111000111111111000000110001111111111100110000001111111100111111100111111111111111111111111000111100000000000000000001111111111",
             "11111111111111001111000000011111011111111111110000000000000001111111111111100001111111110000001100011111111111001100000011111111101111111110011111111111111110111110001111100000000000000000001111111111",
             "11111111111111111100000000000011111111111110000000000000000000000111111000000011111111100000011001111111111110011000000111111111011111111111001111111111101111111000111111110000000000000000011111111111",
             "11111111111111110000111111110001111111111100000100000000000000000000000000110111111111000000110011111111111100110000001111111100110000000000000101110111111111100011111111111000000000000000111111111111",
             "11111111111111100011111111111000111111110000100000000000000000001111111111100111111110000001100111111111111001100000011111111100000001111110000001111111111100000111111111111100000000000011111111111111",
             "11111111111111000111111111111110011111000010000000000000000000000111111111001111111100000011001111111111100011000000111111111000011111111111111000000000000000111111111111101111100000001111011111111111",
             "11111111111111001111111111111110011110001100000000000000000000000011111110111111111000000110011111111111000110000001111111110001111111111111111111000000001111111111111111100011111111111110011111111111",
             "11111111111110011111111111111011001100010000000000000000000000100001111110110001110000001100111111111110001100000011111111100111111111111111111111111111111111111111111111100000111111111000011111111111",
             "11111111111110011111111111111101001110100000000000000000000000010000111111001100011000011000111111111100111000000111111111001111111111111111111111111111111111111111111111100000000000000000011111111111",
             "11111111111110111111111111111001100110000000000000000000000000011000011110111111001000110001111111111001100000001111111100011111111111111111111111111111111111111111111111100000000000000000011111111111",
             "11111111111100111111111111111000100110000000000000000000000000001100001111111111101001100011111111110011000000011111111000111111111111111111111111111111111111111111111111100010000000000000011111111111",
             "11111111111100111111111111111000100110000000000000000000000000000110000111111111101111000111111111100110000000111111110001111111111111111111111111111111111111111111111111100011111100000000011111111111",
             "11111111111100111111111111111000100110000000000000000000000000000011000011111111101110000111111110001100000001111111100011111111111111111111111111111111111111111111111111100011111100000000011111111111",
             "11111111111100111111111111110000100110000000000000000000000000000001100001111111101100001111111100011000000011111111000111111111111111111110000111111111111111111111111111100011111100000000111111111111",
             "11111111111110111111111111110001100110000000000000000000000000000000110000111111011011001111111001110000000111111111001111111111111111111100000001111111111111111111111111100011111100000000111111111111",
             "11111111111110011111111111100001100110000000000000000000000000000000011000011111110111011111110011000000001111111110011111111111111111111000000011101111111111111111111111100011111000000000111111111111",
             "11111111111110011111111110000011001100000000000000000000000000000000001100001111101111011111100110000000011111111100111111111111111111111000000011100001111111111111111111100011111000000000111111111111",
             "11111111111111001111111000000011001100000000000000000000000000000000000110000111111110011111001100000000111111111001111111111111111111110000000111000000011111111111111111000111111000000000111111111111",
             "11111111111111000110000000000110011100000000000000000000000000000000000011000011111110011111001000000001111111110011111111111111111111110000110111000000000011111111111111000111111000000000111111111111",
             "11111111111111100011100000011100111000000000000000000000000000000000000001100001111110011111001000000011111111100111111111111111111111100000111110000000000000111111111111000111111000000001111111111111",
             "11111111111111110001111111110001110000000000000000000000000000000000000000110000111110011111101100000111111111001111111111111111111111100000111110000000000000111111111111000111110000000001111111111111",
             "11111111111111111000001110000011100000000000000000000000000000000000000000011000011110011111100100001111111110011111111111111111111111100000001111001000000001111111111111000111110000000001111111111111",
             "11111111111111111110000000001111000000000000000000000000000000000000000000001100001110011111100110011111111100011111111111111111111111100000000001111111000001111111111111000111110000000001111111111111",
             "11111111111111111111111111111110000000000000000000000000000000000000000000000110000110011111110011111111111100111111111111111111111111110000000000011111000111111111111110001111110000000011111111111111",
             "11111111111111111111111111111000000000000000000000000000000000000000000000000011000010011111111001111111111001111111111111111111111111110000000000000011000011111111111110001111110000000011111111111111",
             "11111111111111111111100100000000000000000000000000000000000000000000000000000000100000011111111100111111110011111111111111111111111100111110000000000000000011111111111110001111100000000011111111111111",
             "11111111111111111111001000000000000000000000000000000000000000000000000000000000010000011111111110011111100111111111111111111111111000011111100000000000000111111111111110001111100000000111111111111111",
             "11111111111111111111001000000000000000000000000000000000000000000000000000000000001000001111111111000111001111111111111111111111110000001111111000000000000111111111111100011111100000000111111111111111",
             "11111111111111111110010000000000000000000000000000000000000000000000000000000000000000001111111111110000011111111111111111111111110000000111111111000000001111111111111100011111000000000111111111111111",
             "11111111111111111110010000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000011111111110000011111111111111100011111000000001111111111111111",
             "11111111111111111110010000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000001111111111111111111111111111000011111000000001111111111111111",
             "11111111111111111100100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000111111111111111111111111111000111110000000001111111111111111",
             "11111111111111111100100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000011111000000011111111111111111111111111000111110000000011111111111111111",
             "11111111111111111100100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000011000000001111111111111111111111110001111100000000011111111111111111",
             "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000111111111111111111111110001111100000000111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000011111111111111111111100001111100000000111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000001111111111111111111100011111000000001111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000111100000000000000000000111111111111111111100011111000000001111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000011110000000000000000000011111111111111111000111110000000011111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000000100111111111111111111111110000000000011111000000000000000000001111111111111111000111110000000011111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000000000111111000000000011111100000000000001111100000001100000000011111111111111110001111100000000111111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000000001111111000000000000111100000011000001111110000000111100000111111111111111110001111000000000111111111111111111111",
             "11111111111111111001000000000000000000000000000000000000000000000000000000000000000001001111111000000000000011100000111000000111111000000011111101111111111111111100011111000000001111111111111111111111",
             "11111111111111111101000000000000000000000000000000000000000000000000000000000000000001001111111000000000000011100000011000000111111100000001111111111111111111111000011110000000011111111111111111111111",
             "11111111111111111100100000000000000000000000000000000000000000000000000000000000000000011111111000001110000011100000011100000111111110000000111111111111111111111000111110000000011111111111111111111111",
             "11111111111111111100100000000000000000000000000000000000000000000000000000000000000010011111111000001110000011110000011100000011111111000000011111111111111111110000111100000000111111111111111111111111",
             "11111111111111111100100000000000000000000000000000000000000000000000000000000000000000111111111000001110000011110000001110000011111111100000011111111111111111110001111000000000111111111111111111111111",
             "11111111111111111100100000000000000000000000000000000000000000000000000000000000000100111111111000001110000011111000001110000001111111110000111111111111111111100001111000000001111111111111111111111111",
             "11111111111111111110110000000000000000000000000000000000000000000000000000000000001001111111111000001110000011111000000110000001111111111001111111111111111111000011110000000011111111111111111111111111",
             "11111111111111111110010000000000000000000000000000000000000000000000000000000000000001111111111000001110000011111000000111000001111111111111111111111111111111000111100000000111111111111111111111111111",
             "11111111111111111110011000000000000000000000000000000000000000000000000000000000010011111111111000001110000011111100000111000000111111111111111111111111111110001111100000000111111111111111111111111111",
             "11111111111111111111001000000000000000000000000000000000000000000000000000000000100111111111111000000000000011111100000011100000111111111111111111111111111100001111000000001111111111111111111111111111",
             "11111111111111111111001000000000000000000000000000000000000000000000000000000001000111111111111000000000000011111110000011100000111111111111111111111111111000011110000000011111111111111111111111111111",
             "11111111111111111111100100000000000000000000000000000000000000000000000000000010001111111111111000000000000111111110000001000000111111111111111111111111110000111100000000111111111111111111111111111111",
             "11111111111111111111100110000000000000000000000000000000000000000000000000000100011111111111111000000000011111111110000000000000111111111111111111111111100001111000000000111111111111111111111111111111",
             "11111111111111111111110010000000000000000000000000000000000000000000000000001000111111111111111000001111111111111111000000000001111111111111111111111111100001110000000001111111111111111111111111111111",
             "11111111111111111111111001000000000000000000000000000000000000000000000000010001111111111111111000001111111111111111000000000111111111111111111111111111000011110000000011111111111111111111111111111111",
             "11111111111111111111111001100000000000000000000000000000000000000000000000100011111111111111111000001111111111111111100000111111111111111111111111111110000111100000000111111111111111111111111111111111",
             "11111111111111111111111100110000000000000000000000000000000000000000000001000111111111111111111000001111111111111111111111111111111111111111111111111100001111000000001111111111111111111111111111111111",
             "11111111111111111111111110010000000000000000000000000000000000000000000010001111111111111111111000001111111111111111111111111111111111111111111111111000011110000000011111111111111111111111111111111111",
             "11111111111111111111111110001000000000000000000000000000000000000000000100011111111111111111111000001111111111111111111111111111111111111111111111110000111100000000111111111111111111111111111111111111",
             "11111111111111111111111111000110000000000000000000000000000000000000001000111111111111111111111111111111111111111111111111111111111111111111111111000001110000000001111111111111111111111111111111111111",
             "11111111111111111111111111100011000000000000000000000000000000000000110001111111111111111111111111111111111111111111111111111111111111111111111110000011100000000011111111111111111111111111111111111111",
             "11111111111111111111111111110001100000000000000000000000000000000001000111111111111111111111111111111111111111111111111111111111111111111111111100000111000000000111111111111111111111111111111111111111",
             "11111111111111111111111111111100011000000000000000000000000000000110001111111111111111111111111111111111111111111111111111111111111111111111111000011110000000011111111111111111111111111111111111111111",
             "11111111111111111111111111111110001100000000000000000000000000011000011111111111111111111111111111111111111111111111111111111111111111111111100000111100000000111111111111111111111111111111111111111111",
             "11111111111111111111111111111111100011000000000000000000000001100001111111111111111111111111111111111111111111111111111111111111111111111111000001110000000001111111111111111111111111111111111111111111",
             "11111111111111111111111111111111110000111000000000000000000110000011111111111111111111111111111111111111111111111111111111111111111111111100000011100000000011111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111100000111100000000011111000011111111111111111111111111111111111111111111111111111111111111111111111111000001110000000001111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111000000111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111100000011100000000011111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000001110000000001111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111000000011000000000011111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001110000000001111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111000000000111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111000000011100000000011111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111000000001100000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111000000000110000000000111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111110000000000110000000000011111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111000000000000100000000000011111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111110000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");  





				 
 label_0 <= (
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
"111111111111111111111111111111111111111001111111111111111111111111111111111111111111", 
"111111111111111111111111111111100000000000000000011111111111111111111111111111111111", 
"111111111111111111111111111100000000000000000000000011111111111111111111111111111111", 
"111111111111111111111111100000000000000000000000000000011111111111111111111111111111", 
"111111111111111111111110000000000000000000000000000000000111111111111111111111111111", 
"111111111111111111111100000000000000000000000000000000000011111111111111111111111111", 
"111111111111111111111000000000000000000000000000000000000000111111111111111111111111", 
"111111111111111111100000000000000000000000000000000000000000011111111111111111111111", 
"111111111111111111000000000000000000000000000000000000000000001111111111111111111111", 
"111111111111111111000000000000000000000000000000000000000000000111111111111111111111", 
"111111111111111110000000000000000000000000000000000000000000000011111111111111111111", 
"111111111111111100000000000000000000000000000000000000000000000001111111111111111111", 
"111111111111111100000000000000000000000000000000000000000000000001111111111111111111", 
"111111111111111000000000000000000000000000000000000000000000000000111111111111111111", 
"111111111111111000000000000000000000000000000000000000000000000000111111111111111111", 
"111111111111110000000000000000000000000000000000000000000000000000011111111111111111", 
"111111111111110000000000000000000000000000000000000000000000000000011111111111111111", 
"111111111111110000000000000000000000000111000000000000000000000000011111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111100000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111100000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111110000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111100000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111100000000000000000000000000111111111111111", 
"111111111111000000000000000000000000001111100000000000000000000000000111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
"111111111111110000000000000000000000000111000000000000000000000000001111111111111111", 
"111111111111110000000000000000000000000000000000000000000000000000011111111111111111", 
"111111111111110000000000000000000000000000000000000000000000000000011111111111111111", 
"111111111111111000000000000000000000000000000000000000000000000000011111111111111111", 
"111111111111111000000000000000000000000000000000000000000000000000111111111111111111", 
"111111111111111100000000000000000000000000000000000000000000000000111111111111111111", 
"111111111111111100000000000000000000000000000000000000000000000001111111111111111111", 
"111111111111111110000000000000000000000000000000000000000000000011111111111111111111", 
"111111111111111111000000000000000000000000000000000000000000000011111111111111111111", 
"111111111111111111000000000000000000000000000000000000000000000111111111111111111111", 
"111111111111111111100000000000000000000000000000000000000000001111111111111111111111", 
"111111111111111111110000000000000000000000000000000000000000011111111111111111111111", 
"111111111111111111111100000000000000000000000000000000000000111111111111111111111111", 
"111111111111111111111110000000000000000000000000000000000011111111111111111111111111", 
"111111111111111111111111100000000000000000000000000000000111111111111111111111111111", 
"111111111111111111111111111000000000000000000000000000111111111111111111111111111111", 
"111111111111111111111111111111000000000000000000000111111111111111111111111111111111", 
"111111111111111111111111111111111111000000000111111111111111111111111111111111111111", 
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111"); 
 
label_1 <= (
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111000000000000000011111111111111111111111111111",
"111111111111111111111111111111111111110000000000000000011111111111111111111111111111",
"111111111111111111111111111111111111100000000000000000011111111111111111111111111111",
"111111111111111111111111111111111111000000000000000000011111111111111111111111111111",
"111111111111111111111111111111111110000000000000000000011111111111111111111111111111",
"111111111111111111111111111111111100000000000000000000011111111111111111111111111111",
"111111111111111111111111111111111000000000000000000000011111111111111111111111111111",
"111111111111111111111111111111100000000000000000000000011111111111111111111111111111",
"111111111111111111111111111111000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111100000000000000000000000000011111111111111111111111111111",
"111111111111111111111111110000000000000000000000000000011111111111111111111111111111",
"111111111111111111111111000000000000000000000000000000011111111111111111111111111111",
"111111111111111111111100000000000000000000000000000000011111111111111111111111111111",
"111111111111111111100000000000000000000000000000000000011111111111111111111111111111",
"111111111111111100000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111100000000000000000000000000000000000000000011111111111111111111111111111",
"111111111111111111111111000000000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111000000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111100000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111100000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
		

label_2 <= (
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111011111111111111111111111111111111111111111111111",
"111111111111111111111111111100000000000000000011111111111111111111111111111111111111",
"111111111111111111111111100000000000000000000000001111111111111111111111111111111111",
"111111111111111111111110000000000000000000000000000011111111111111111111111111111111",
"111111111111111111111000000000000000000000000000000000111111111111111111111111111111",
"111111111111111111110000000000000000000000000000000000001111111111111111111111111111",
"111111111111111111100000000000000000000000000000000000000111111111111111111111111111",
"111111111111111111000000000000000000000000000000000000000011111111111111111111111111",
"111111111111111110000000000000000000000000000000000000000001111111111111111111111111",
"111111111111111100000000000000000000000000000000000000000000111111111111111111111111",
"111111111111111000000000000000000000000000000000000000000000011111111111111111111111",
"111111111111110000000000000000000000000000000000000000000000001111111111111111111111",
"111111111111110000000000000000000000000000000000000000000000001111111111111111111111",
"111111111111100000000000000000000000000000000000000000000000000111111111111111111111",
"111111111111100000000000000000000000000000000000000000000000000111111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111111000000000000000000000000111000000000000000000000000011111111111111111111",
"111111111110000000000000000000000001111110000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111111000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111111000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000000111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000000111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000000111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000000111111111111111111",
"111111111110000000000000000000000011111110000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111100000000000000000000000001111111111111111111",
"111111111110000000000000000000000011111100000000000000000000000001111111111111111111",
"111111111100000000000000000000000011111100000000000000000000000001111111111111111111",
"111111111100000000000000000000000011111000000000000000000000000001111111111111111111",
"111111111100000000000000000000000011111000000000000000000000000001111111111111111111",
"111111111100000000000000000000000011110000000000000000000000000001111111111111111111",
"111111111100000000000000000000000011110000000000000000000000000011111111111111111111",
"111111111111111111111111111111111111100000000000000000000000000011111111111111111111",
"111111111111111111111111111111111111100000000000000000000000000011111111111111111111",
"111111111111111111111111111111111111000000000000000000000000000111111111111111111111",
"111111111111111111111111111111111111000000000000000000000000000111111111111111111111",
"111111111111111111111111111111111110000000000000000000000000000111111111111111111111",
"111111111111111111111111111111111110000000000000000000000000001111111111111111111111",
"111111111111111111111111111111111100000000000000000000000000001111111111111111111111",
"111111111111111111111111111111111100000000000000000000000000011111111111111111111111",
"111111111111111111111111111111111000000000000000000000000000011111111111111111111111",
"111111111111111111111111111111111000000000000000000000000000111111111111111111111111",
"111111111111111111111111111111110000000000000000000000000000111111111111111111111111",
"111111111111111111111111111111100000000000000000000000000001111111111111111111111111",
"111111111111111111111111111111100000000000000000000000000001111111111111111111111111",
"111111111111111111111111111111000000000000000000000000000011111111111111111111111111",
"111111111111111111111111111111000000000000000000000000000111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000000111111111111111111111111111",
"111111111111111111111111111110000000000000000000000000001111111111111111111111111111",
"111111111111111111111111111100000000000000000000000000001111111111111111111111111111",
"111111111111111111111111111000000000000000000000000000011111111111111111111111111111",
"111111111111111111111111111000000000000000000000000000111111111111111111111111111111",
"111111111111111111111111110000000000000000000000000000111111111111111111111111111111",
"111111111111111111111111100000000000000000000000000001111111111111111111111111111111",
"111111111111111111111111100000000000000000000000000011111111111111111111111111111111",
"111111111111111111111111000000000000000000000000000011111111111111111111111111111111",
"111111111111111111111111000000000000000000000000000111111111111111111111111111111111",
"111111111111111111111110000000000000000000000000001111111111111111111111111111111111",
"111111111111111111111110000000000000000000000000001111111111111111111111111111111111",
"111111111111111111111100000000000000000000000000011111111111111111111111111111111111",
"111111111111111111111000000000000000000000000000111111111111111111111111111111111111",	
"111111111111111111111000000000000000000000000000111111111111111111111111111111111111",
"111111111111111111110000000000000000000000000001111111111111111111111111111111111111",
"111111111111111111110000000000000000000000000011111111111111111111111111111111111111",
"111111111111111111100000000000000000000000000011111111111111111111111111111111111111",
"111111111111111111000000000000000000000000000111111111111111111111111111111111111111",
"111111111111111111000000000000000000000000001111111111111111111111111111111111111111",
"111111111111111110000000000000000000000000001111111111111111111111111111111111111111",
"111111111111111100000000000000000000000000011111111111111111111111111111111111111111",
"111111111111111100000000000000000000000000111111111111111111111111111111111111111111",
"111111111111111000000000000000000000000000111111111111111111111111111111111111111111",
"111111111111111000000000000000000000000001111111111111111111111111111111111111111111",
"111111111111110000000000000000000000000011111111111111111111111111111111111111111111",
"111111111111100000000000000000000000000111111111111111111111111111111111111111111111",
"111111111111100000000000000000000000000111111111111111111111111111111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111110000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111100000000000000000000000000000000000000000000000000000011111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

label_3 <= (
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111110000000111111111111111111111111111111111111111111",
"111111111111111111111111111000000000000000000000011111111111111111111111111111111111",
"111111111111111111111110000000000000000000000000000001111111111111111111111111111111",
"111111111111111111111000000000000000000000000000000000011111111111111111111111111111",
"111111111111111111100000000000000000000000000000000000000111111111111111111111111111",
"111111111111111110000000000000000000000000000000000000000001111111111111111111111111",
"111111111111111100000000000000000000000000000000000000000000111111111111111111111111",
"111111111111111000000000000000000000000000000000000000000000011111111111111111111111",
"111111111111111000000000000000000000000000000000000000000000001111111111111111111111",
"111111111111110000000000000000000000000000000000000000000000001111111111111111111111",
"111111111111110000000000000000000000000000000000000000000000000111111111111111111111",
"111111111111100000000000000000000000000000000000000000000000000011111111111111111111",
"111111111111100000000000000000000000000000000000000000000000000011111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000001111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000001111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000001111111111111111111",
"111111111111000000000000000000000000000000000000000000000000000000111111111111111111",
"111111111110000000000000000000000000001110000000000000000000000000111111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000111111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000111111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000111111111111111111",
"111111111111111111111111111111111111111111000000000000000000000000111111111111111111",
"111111111111111111111111111111111111111111000000000000000000000000111111111111111111",
"111111111111111111111111111111111111111110000000000000000000000000111111111111111111",
"111111111111111111111111111111111111111110000000000000000000000001111111111111111111",
"111111111111111111111111111111111111100000000000000000000000000001111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000011111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000111111111111111111111",
"111111111111111111111111111100000000000000000000000000000000001111111111111111111111",
"111111111111111111111111111100000000000000000000000000000000011111111111111111111111",
"111111111111111111111111111100000000000000000000000000000001111111111111111111111111",
"111111111111111111111111111100000000000000000000000000000011111111111111111111111111",
"111111111111111111111111111100000000000000000000000000000000011111111111111111111111",
"111111111111111111111111111100000000000000000000000000000000001111111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000111111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000011111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000001111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000001111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000000111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000000111111111111111111",
"111111111111111111111111111100000000000000000000000000000000000000111111111111111111",
"111111111111111111111111111110000000000000000000000000000000000000011111111111111111",
"111111111111111111111111111111111111111000000000000000000000000000011111111111111111",
"111111111111111111111111111111111111111100000000000000000000000000011111111111111111",
"111111111111111111111111111111111111111110000000000000000000000000011111111111111111",
"111111111111111111111111111111111111111110000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000011111111111111111",
"111111111110000000000000000000000000011111000000000000000000000000001111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",		
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000001111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",	
"111111111110000000000000000000000000111111000000000000000000000000011111111111111111",	
"111111111111000000000000000000000000011111000000000000000000000000011111111111111111",	
"111111111111000000000000000000000000011111000000000000000000000000011111111111111111",	
"111111111111000000000000000000000000011111000000000000000000000000011111111111111111",	
"111111111111000000000000000000000000011110000000000000000000000000111111111111111111",	
"111111111111000000000000000000000000000000000000000000000000000000111111111111111111",	
"111111111111100000000000000000000000000000000000000000000000000000111111111111111111",	
"111111111111100000000000000000000000000000000000000000000000000000111111111111111111",	
"111111111111100000000000000000000000000000000000000000000000000001111111111111111111",	
"111111111111110000000000000000000000000000000000000000000000000001111111111111111111",	
"111111111111110000000000000000000000000000000000000000000000000011111111111111111111",	
"111111111111111000000000000000000000000000000000000000000000000011111111111111111111",	
"111111111111111000000000000000000000000000000000000000000000000111111111111111111111",	
"111111111111111100000000000000000000000000000000000000000000001111111111111111111111",	
"111111111111111110000000000000000000000000000000000000000000011111111111111111111111",	
"111111111111111111000000000000000000000000000000000000000000111111111111111111111111",	
"111111111111111111110000000000000000000000000000000000000001111111111111111111111111",	
"111111111111111111111000000000000000000000000000000000000011111111111111111111111111",	
"111111111111111111111110000000000000000000000000000000001111111111111111111111111111",	
"111111111111111111111111100000000000000000000000000000111111111111111111111111111111",	
"111111111111111111111111111100000000000000000000001111111111111111111111111111111111",	
"111111111111111111111111111111111100000000000111111111111111111111111111111111111111",	
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",	
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111",	
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111");					 

StartGameLabel <=("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111100111111111111111111111111001111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111100000011111000011111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111100111111111111111111111100001111111111111111111110110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111110001111100011110011111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111100111111111111111111111111001111111111111111111101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111100111111110011110011111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111001111111111011110011111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111011111111111111111001111111111111111111001111111111111111111111111111111111111111111111011111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111110001111111111111110011111111111111111111111111111111111111111111111111111111111111111111101111110011111111111111111111111111111111111111111111111111111111111111111110011111111111111111001111111111111111111001111111111111111111111111111111111111111111110011111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111110011111111111101110011111111111111111111111111111111111111111111111111111111111111111111001111110011111111111111111111111111111111111111111111111111111111111111111100011111111111111111001111111111111111111001111111111111111111111111111111111111111111110011111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111100011111111111111110011100011111100000111111001110001111111100001111111110000111111111110000001110011000011111110000111111111111100000011000001100000111000011100111000000011110000011111001110001111111111100000001111100000111111001100111111111110000011000000011110000011111101100010000001111111111100000111111110000011111100110000111000011111110000011111111111111111111111111",
					   "1111111111111111111111111100011111111111111110010010001111001110011110001000000111110011100000111001110001111111111101111110010100011111001110001111111111001110011100011110001111100110000111110011111101110001111001001000111111111111001111110011110011100001000011111111001110011110011111001110001110001000011001111111111111001110000011001110001110000101000110000001111101110001111111111111111111111111",
					   "1111111111111111111111111100011111111111111110001111001111001111001111000111100111100011110011110011111001111111111101111110011111001111011111001111111111011111011110011111001111101111100111110011111011111001111000111100111111111111001111110111111001111000110111111111011111011110011111001111001111000111111001111111111110011111001111001111001111000111110001111001111011111000111111111111111111111111",
					   "1111111111111111111111111100011111111111111110011111001111011111001111001111100111100111110011110111111000111111111101111110011111001110011111000111111111011111011110011111001111101111100111110011110011111001111001111100111111111111001111100111111000111001111111111111001111111110011111001111001111000111111001111111111110011111001111001111001111100111110011111001110011111000111111111111111111111111",
					   "1111111111111111111111111100011111111111111110011111001111111100001111001111100111100111110011110000000000111111111101111110011111001110000000000111111111000111111111001111000111011111100111110011110011111111111001111100111111111111001111100111111000111001111111111111000111111110011111111110001111001111111001111111111110011111001111111110001111100111110011111001110000000000111111111111111111111111",
					   "1111111111111111111111111100011111111111111110011111001111110011001111001111100111100011110011110111111111111111111101111110011111001110011111111111111111100001111111001110100111011111100111110011110011111111111001111100111111111111001111100111111100111001111111111111100001111110011111110001001111001111111001111111111110011111001111110001001111100111110011111001110011111111111111111111111111111111",
					   "1111111111111111111111111110011111111111111110011111001111001111001111001111100111110011100011110011111111111111111101111110011111001110011111111111111111111000011111000110110011011111100111110011110011111111111001111100111111111111001111100111111100111001111111111111111000011110011111100111001111001111111001111111111111001110011111100111001111100111110011111001110011111111111111111111111111111111",
					   "1111111111111111111111111110001111111111111110011111001110011111001111001111100111111000001111110011111111111111111101111110011111001110011111111111111111111110011111100101110010111111100111110011110011111111111001111100111111111111001111100111111100111001111111111111111110001110011111001111001111001111111001111111111111100000111111001111001111100111110011111001110011111111111111111111111111111111",
					   "1111111111111111111111111111001111111111011110011111001110011111001111001111100111110111111111110001111111111111111101111110011111001110001111110111111111111111001111100001110000111111100111110011110001111111111001111100111111111111001111100111111001111001111111111111111111001110011110011111001111001111111001111111111111011111111110011111001111100111110011111001110001111110111111111111111111111111",
					   "1111111111111111111111111111000011111110011110011111001110011110001111001111100111100111111111110000111001111111111100111110011111001111000011001111111111011111001111110011111001111111100111110011111000111101111001111100111111111111001111100011111001111001111111111111011111001110011110001111001111001111111001111111111110011111111110001111001111100111110011111001111000011101111111111111111111111111",
					   "1111111111111111111111111111110000111101111110011111000110000001000111000111100011100000000011111000000011111111111100001100011111001111000000011111111111001110011111110011111001111111000111110000111000000011111001111100011111111111000111110001110011111000111111111111001111011110000011000101000011000111111000101111111110000000001111000101000011000111110011111000111100000001111111111111111111111111",
					   "1111111111111111111111111111111100000011111000000100000011000011001100000011000001110000000000111110000111111111111100011000000100000011110000111111111111000000111111111111111111111110000001111001111110000111100000010000001111111100000001111100001111100000011111111111000000111111000111000011000100000011111100011111111111000000000111000011000110000001000000100000011110000111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111011111011111011111011111011111011111011111011111011001011111010111011111011111111111111101111101111101111101111101111111111111101111101111101111101111101111101111101111101111101111101111101111111111111111011111011111011111011111011111111111001111001111001111001111001111001111001111111111100111011110011111011111011111011111011111011111011111011111111111111111111111111",
					   "1111111111111111111111111111111101111101111101111101111101111101111101111101111101000101111101111101111101111111111111110111110111110111110111110111111111111110111110111110111110111110111110111110111110111110111110111110111011111111111101111101111101111101111101111100110010110010110010110010110010110010110010111011111100111101100101111101111101111101111101111101111101111101110111111111111111111111",
					   "1111111111111111111111111101101111101111101111101111101111101111101111101111101111100000000001101111101110111111110110111110111110111110111110111011111110110111110111110111110111110111110111110111110111110111110111110111110111111101101111101111101111101111101110111110110110010110010110010110010110010110010110010111111100000000001111101111101111101111101111101111101111101111101111111111111111111111",
					   "1111111111111111111111111111011111011111011111011111011111011111011111011111011111010000001111011111011111111111111101111101111101111101111101111111111111101111101111101111101111101111101111101111101111101111101111101111101111111111011111011111011111011111011111111111001111001111001111001111001111001111001111001111111110000000011111011111011111011111011111011111011111011111011111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
					   "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
					   
P1_Won_Label <= (
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1100000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111",
"1100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111",
"1100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111",
"1110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111",
"1111000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111",
"1111000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111000000000000000111111",
"1111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000000000000000000000000000000000000000000000001111110000000000000000001111111111111111111111111111111111111111111111100000000000000000001111111111111111111000000000000000000000011111111110000000000000000000000100000000000000000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000000111111111111111111111100000000000000000001111110000000000000000001111111111111111111111111111111111111111111111000000000000000000001111111111111111110000000000000000000000011111111110000000000000000000000100000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111100000000000000001111110000000000000000001111111111111111111111111111111111111111111111000000000000000000001111111111111111110000000000000000000000011111111110000000000000000000000100000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111110000000000000000111111000000000000000111111111111111111111111111111111111111111111111100000000000000000011111111111111111111100000000000000000000111111111111100000000000000000011111000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111111000000000000000111111100000000000001111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111000000000000000011111111111111110000000000000001111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111111000000000000000111111100000000000001111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111100000000000000011111111111111110000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111111100000000000000111111100000000000001111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111110000000000000001111111111111100000000000000111111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111111100000000000000111111100000000000001111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111000000000000001111111111111000000000000000111111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111111100000000000000111111100000000000001111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111000000000000000111111111111000000000000001111111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111110000000000000000000000111111",
"1111000000000000001111111111111111111111111111100000000000000111111100000000000001111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000000000111111111110000000000000011111111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000011110000000000000111111",
"1111000000000000001111111111111111111111111111000000000000000111111100000000000001111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111110000000000000011111111100000000000000111111111111100000000000001111111111111111111111111110000011111111100000000000000111111111111111110000000000000000001111111111111111111111111111111111111111110000111110000000000000111111",
"1111000000000000001111111111111111111111111111000000000000000111111100000000000001111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111110000000000000001111111100000000000000111111111111100000000000001111111111111111111111111111100011111111100000000000001111111111111111111111000000000000001111111111111111111111111111111111111111110000111110000000000000111111",
"1111000000000000001111111111111111111111111110000000000000001111111100000000000001111111111111111111111111111111111111111111111111000000000000000000000111111111111111111111111111000000000000000111111000000000000001111111111111100000000000001111111111111111111111111111100011111111100000000000001111111111111111111111100000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111100000000000000001111111100000000000001111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111100000000000000111110000000000000011111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111111111111111100000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000111000000000000000000000001111111100000000000001111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111110000000000000011110000000000000111111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111111111111111100000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000000011111111100000000000001111111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111110000000000000001100000000000000111111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111111111111111100000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000000111111111100000000000001111111111111111111111111111111111111111111111100000000000100000000000001111111111111111111111111111000000000000000000000000000001111111111111111100000000000001111111111111111111001111111111111111111100000000000001111111111111111111111100000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000000111111111100000000000001111111111111111111111111111111111111111111111000000000000110000000000000111111111111111111111111111100000000000000000000000000011111111111111111100000000000001111111111111111110001111111111111111111100000000000001111111111111111111111100000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000001111111111100000000000001111111111111111111111111111111111111111111111000000000001110000000000000111111111111111111111111111110000000000000000000000000011111111111111111100000000000001111111111111111110001111111111111111111100000000000001111111111111111111110000000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000011111111111100000000000001111111111111111111111111111111111111111111110000000000001111000000000000011111111111111111111111111110000000000000000000000000111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000000111111111111100000000000001111111111111111111111111111111111111111111110000000000011111000000000000011111111111111111111111111111000000000000000000000001111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000001111111111111100000000000001111111111111111111111111111111111111111111100000000000011111100000000000001111111111111111111111111111100000000000000000000011111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000000011111111111111100000000000001111111111111111111111111111111111111111111100000000000111111100000000000001111111111111111111111111111100000000000000000000011111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000000001111111111111111100000000000001111111111111111111111111111111111111111111000000000000111111110000000000000111111111111111111111111111110000000000000000000111111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000000000000001111111111111111111100000000000001111111111111111111111111111111111111111111000000000001111111110000000000000111111111111111111111111111111000000000000000001111111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000000000000000000000111111111111111111111111111111100000000000001111111111111111111111111111111111111111110000000000001111111111000000000000011111111111111111111111111111100000000000000011111111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111110000000000011111111111000000000000011111111111111111111111111111100000000000000011111111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111100000000000011111111111100000000000001111111111111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111100000000000011111111111100000000000001111111111111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000001111111111111111111100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111110001111111111111111111100000000000000111111111000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111001111111111111111111100000000000001111111111100000000000000111111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111100000000000000111111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111110000000000000011111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111111000000000000001111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111111100000000000000111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111111111111111111111111100000000000001111111111111100000000000000111111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111001111111000000000000000000000000000000000000000000000111111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111111111111110001111111100000000000001111111111111110000000000000011111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000001111111111111111111111111110001111110000000000001111111111111111111110000000000000011111111111111111111111110000000000000111111111111111111111111100000000000001111111111111111111111111111110001111111100000000000001111111111111111000000000000001111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001111110000000000001111111111111111111111000000000000011111111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000001111111100000000000001111111111111111000000000000001111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001111100000000000011111111111111111111111000000000000001111111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000001111111100000000000001111111111111111100000000000000111111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001111100000000000011111111111111111111111100000000000000111111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000001111111100000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001111000000000000111111111111111111111111100000000000000111111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000001111111100000000000001111111111111111111000000000000001111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001111000000000000111111111111111111111111110000000000000011111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000001111111100000000000001111111111111111111000000000000000111111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001110000000000000111111111111111111111111110000000000000011111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000001111111100000000000001111111111111111111100000000000000011111111111111111111111111111111111111111111111111110000000000000111111",
"1111000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001110000000000000111111111111111111111111110000000000000001111111111111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000001111111100000000000001111111111111111111100000000000000001111111111111111111111111111111111111111111111111100000000000000011111",
"1100000000000000000011111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000011111111111111111100000000000000011111111111111111111110000000000000000000000000000000000000000000000001111111000000000000000011111111111111111000000000000000000011111111111111111111111111111111111111111111111000000000000000001111",
"1100000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111110000000000000000000111111111111111111100000000000000000000000000000000000000000000000001111110000000000000000001111111111111110000000000000000000001111111111111111111111111111111111111111111110000000000000000000111",
"1100000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111110000000000000000000111111111111111111100000000000000000000000000000000000000000000000001111110000000000000000001111111111111110000000000000000000001111111111111111111111111111111111111111111110000000000000000000111",
"1100000000000000000011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111000000000000000001111111111111111111110000000000000000000000000000000000111111111000001111110000000000000000011111111111111111000000000000000000001111111111111111111111111111111111111111111111000000000000000000111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111110000000000000000000011111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111110000000000000000000011111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111100000000000000000000011111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111000000000000000000111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111000000000000000001111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111000000000000000001111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111000000000000000001111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111110000000000000000001111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111110000000000000000000111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111110000000000000000000111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111110000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111100000000000000000000011111111111111111110000000000000011111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111100000000000000000000011111111111111111110000000000000011111111111111111111111000000000000000000000011111111111111111111111000000000000000000011111111111111111111000000000000000001111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111100000000000000000000011111111111111111100000000000000111111111111111111111100000000000000000000000000111111111111111111111000000000000000000011111111111111111111000000000000000001111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111000000000000000000000001111111111111111100000000000000111111111111111111110000000000000000000000000000001111111111111111111000000000000000000011111111111111111111100000000000000001111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111000000000000000000000001111111111111111000000000000001111111111111111111000000000000000000000000000000000111111111111111111110000000000000001111111111111111111111110000000000000111111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110000000000000001111111111111110000000000000000000000001111111111111111000000000000001111111111111111100000000000000000000000000000000000001111111111111111110000000000000000111111111111111111111111000000000000111111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110000000000000001111111111111110000000000000000000000000111111111111111000000000000001111111111111111000000000000000000000000000000000000000111111111111111110000000000000000011111111111111111111111000000000000111111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111000000000000001111111111111110000000000000000000000000111111111111110000000000000011111111111111110000000000000000000000000000000000000000011111111111111110000000000000000001111111111111111111111000000000000111111111111111111111111111111111111100000000000111111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111000000000000000111111111111100000000000000000000000000011111111111110000000000000011111111111111100000000000000000000000000000000000000000001111111111111110000000000000000000111111111111111111111000000000000111111111111111111111111111111111111100000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111100000000000000111111111111100000000000000000000000000011111111111110000000000000011111111111111000000000000000000000000000000000000000000000011111111111110000000000000000000011111111111111111111000000000000111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111100000000000000111111111111000000000000001000000000000011111111111100000000000000111111111111110000000000000000000001111110000000000000000000011111111111110000000000000000000001111111111111111111000000000000111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111100000000000000011111111111000000000000011000000000000001111111111100000000000000111111111111110000000000000000001111111111111000000000000000001111111111110000000000000000000000111111111111111111000000000000111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111110000000000000011111111111000000000000011000000000000001111111111100000000000001111111111111100000000000000000111111111111111100000000000000000111111111110000000000000000000000011111111111111111000000000000111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111110000000000000011111111110000000000000111100000000000001111111111000000000000001111111111111100000000000000011111111111111111111000000000000000011111111110000000000000000000000011111111111111111000000000000111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111000000000000001111111110000000000000111100000000000000111111111000000000000001111111111111000000000000000111111111111111111111100000000000000011111111110000000000000000000000001111111111111111000000000000111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111000000000000001111111110000000000000111100000000000000111111110000000000000011111111111111000000000000001111111111111111111111110000000000000011111111110000000000000000000000000111111111111111000000000000111111111111111111111111111111111111110000000001111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111000000000000001111111100000000000001111110000000000000111111110000000000000011111111111110000000000000011111111111111111111111111000000000000001111111110000000000000000000000000011111111111111000000000000111111111111111111111111111111111111110000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111100000000000000111111100000000000001111110000000000000011111110000000000000111111111111110000000000000011111111111111111111111111000000000000001111111110000000000000000000000000001111111111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111100000000000000111111000000000000001111111000000000000011111100000000000000111111111111110000000000000111111111111111111111111111100000000000001111111110000000000000000000000000000111111111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111100000000000000011111000000000000011111111000000000000001111100000000000000111111111111110000000000000111111111111111111111111111100000000000000111111110000000000001000000000000000011111111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111110000000000000011111000000000000011111111000000000000001111100000000000001111111111111100000000000000111111111111111111111111111110000000000000111111110000000000001100000000000000001111111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111110000000000000011110000000000000111111111100000000000001111000000000000001111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001110000000000000000111111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111000000000000001110000000000000111111111100000000000000111000000000000011111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001111000000000000000011111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111000000000000001100000000000000111111111100000000000000111000000000000011111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001111100000000000000001111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111000000000000001100000000000001111111111110000000000000110000000000000011111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001111110000000000000000111111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111100000000000000100000000000001111111111110000000000000010000000000000111111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001111111000000000000000011111000000000000111111111111111111111111111111111111111000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111000000000000000000000000000111111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001111111100000000000000001111000000000000111111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111000000000000000000000000000111111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001111111110000000000000000111000000000000111111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111000000000000000000000000001111111111111111100000000000001111111111111111111111111111110000000000000111111110000000000001111111111000000000000000011000000000000111111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000111111111111111111111111111110000000000000111111110000000000001111111111100000000000000001000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111110000000000000111111111111111111111111111100000000000000111111110000000000001111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111110000000000000011111111111111111111111111100000000000000111111110000000000001111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111110000000000000011111111111111111111111111000000000000001111111110000000000001111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111110000000000000001111111111111111111111111000000000000001111111110000000000001111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111000000000000000000000111111111111111111111000000000000000111111111111111111111110000000000000001111111110000000000001111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111000000000000000000001111111111111111111111000000000000000111111111111111111111100000000000000011111111110000000000001111111111111111100000000000000000000000111111111111111111111111111111111111111100000001111111111111111111111111000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111000000000000000000001111111111111111111111100000000000000001111111111111111111000000000000000011111111110000000000001111111111111111110000000000000000000000111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111100000000000000000001111111111111111111111100000000000000000111111111111111100000000000000000111111111110000000000001111111111111111111000000000000000000000111111111111111111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111100000000000000000011111111111111111111111110000000000000000001111111111110000000000000000001111111111110000000000001111111111111111111000000000000000000000111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000001111111111110000000000001111111111111111111100000000000000000000111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111110000000000000000111111111111111111111111111100000000000000000000000000000000000000000000011111111111110000000000001111111111111111111110000000000000000000111111111111111111111111111111111110000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111110000000000000000111111111111111111111111111110000000000000000000000000000000000000000000111111111111110000000000001111111111111111111111000000000000000000111111111111111111111111111111111110000000000000001111111111111111100000000000000001111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111000000000000000111111111111111111111111111111000000000000000000000000000000000000000001111111111111110000000000001111111111111111111111100000000000000000111111111111111111111111111111111110000000000000001111111111111111100000000000000001111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111000000000000001111111111111111111111111111111110000000000000000000000000000000000000011111111111111110000000000001111111111111111111111110000000000000000111111111111111111111111111111111110000000000000001111111111111111100000000000000001111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111000000000000001111111111111111111111111111111111000000000000000000000000000000000000111111111111111110000000000001111111111111111111111111000000000000000111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111110000000000000000111111111111111111111111111111111100000000000000000000000000000000011111111111111111110000000000000111111111111111111111111100000000000000111111111111111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111000000000000000000001111111111111111111111111111111111000000000000000000000000000001111111111111111111000000000000000001111111111111111111110000000000000000001111111111111111111111111111111111000000000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111000000000000000000001111111111111111111111111111111111110000000000000000000000000111111111111111111111000000000000000001111111111111111111110000000000000000001111111111111111111111111111111111100000000000111111111111111111111000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111000000000000000000001111111111111111111111111111111111111110000000000000000000011111111111111111111111000000000000000001111111111111111111110000000000000000001111111111111111111111111111111111110000000001111111111111111111111110000000011111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111000001111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
	

P2_Won_Label <= (
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111111111111111111",
"1110000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111",
"1110000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111",
"1110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111",
"1111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111",
"1111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111",
"1111110000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000001111111111111",
"1111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111",
"1111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111",
"1111110000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000001111111111",
"1111110000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111",
"1111110000000000000000000000000000000000000000000000000000011111000000000000000001111111111111111111111111111111111111111111110000000000000000001111111111111111110000000000000000000001111111111000000000000000000000100000000000000000000000000000000000000000000001111110000000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000111111111100000000000000001111111111",
"1111110000000000000111111111111111111111111000000000000000011111000000000000000001111111111111111111111111111111111111111111110000000000000000001111111111111111110000000000000000000001111111111000000000000000000000100000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000111111111111110000000000000000111111111",
"1111110000000000000111111111111111111111111110000000000000011111100000000000000001111111111111111111111111111111111111111111110000000000000000001111111111111111111000000000000000000001111111111100000000000000000001110000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000011111111111111111100000000000000111111111",
"1111110000000000000111111111111111111111111110000000000000001111110000000000000111111111111111111111111111111111111111111111111100000000000000011111111111111111111110000000000000000111111111111110000000000000000111111000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000001111111111111111111111111111111111000000000001111111111111111111100000000000000111111111",
"1111110000000000000111111111111111111111111111000000000000001111111000000000000111111111111111111111111111111111111111111111111100000000000000111111111111111111111111000000000000000111111111111110000000000000011111111000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000111111111111111111111111111111111100000000011111111111111111111110000000000000111111111",
"1111110000000000000111111111111111111111111111000000000000001111111000000000000111111111111111111111111111111111111111111111111100000000000000111111111111111111111111100000000000000111111111111110000000000000011111111000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000011111111111111111111111111111111110000000111111111111111111111110000000000000111111111",
"1111110000000000000111111111111111111111111111000000000000001111111000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111110000000000000011111111111100000000000000111111111000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000011111111111111111111111111111111111000000111111111111111111111110000000000000111111111",
"1111110000000000000111111111111111111111111111000000000000001111111000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111110000000000000011111111111100000000000001111111111000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000001111111111111111111111111111111111000001111111111111111111111110000000000000111111111",
"1111110000000000000111111111111111111111111111000000000000001111111000000000000111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111000000000000001111111111000000000000011111111111000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000001111111111111111111111111111111111100000111111111111111111111100000000000000111111111",
"1111110000000000000111111111111111111111111111000000000000001111111000000000000111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111100000000000000111111110000000000000011111111111000000000000011111111111111111111111111100001111111100000000000001111111111111111100000000000000000111111111111111111111111111111111110000111111111111111111111100000000000000111111111",
"1111110000000000000111111111111111111111111110000000000000011111111000000000000111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111110000000000000111111110000000000000111111111111000000000000011111111111111111111111111110001111111100000000000011111111111111111111100000000000000111111111111111111111111111111111111000111111111111111111111100000000000000111111111",
"1111110000000000000111111111111111111111111100000000000000011111111000000000000111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111110000000000000011111100000000000001111111111111000000000000011111111111111111111111111110011111111100000000000011111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111000000000000000111111111",
"1111110000000000000111111111111111111111111000000000000000011111111000000000000111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111000000000000001111000000000000011111111111111000000000000011111111111111111111111111111111111111100000000000011111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111110000000000000000111111111",
"1111110000000000000000000000000000000000000000000000000000111111111000000000000111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111100000000000000111000000000000011111111111111000000000000011111111111111111111111111111111111111100000000000011111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111000000000000000001111111111",
"1111110000000000000000000000000000000000000000000000000000111111111000000000000111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111110000000000000110000000000000111111111111111000000000000011111111111111111111111111111111111111100000000000011111111111111111111110000000000000111111111111111111111111111111111111111111111111111111110000000000000000001111111111",
"1111110000000000000000000000000000000000000000000000000001111111111000000000000111111111111111111111111111111111111111111110000000000010000000000001111111111111111111111111110000000000000000000000000001111111111111111000000000000011111111111111111100111111111111111111100000000000011111111111111111111110000000000000111111111111111111111111111111111111111111111111111111000000000000000000011111111111",
"1111110000000000000000000000000000000000000000000000000011111111111000000000000111111111111111111111111111111111111111111100000000000111000000000000111111111111111111111111111000000000000000000000000011111111111111111000000000000011111111111111111000111111111111111111100000000000011111111111111111111100000000000000111111111111111111111111111111111111111111111111111100000000000000000000011111111111",
"1111110000000000000000000000000000000000000000000000000011111111111000000000000111111111111111111111111111111111111111111100000000000111000000000000011111111111111111111111111100000000000000000000000011111111111111111000000000000000000000000000000000111111111111111111100000000000001111111111111111110000000000000001111111111111111111111111111111111111111111111111100000000000000000000000111111111111",
"1111110000000000000000000000000000000000000000000000000111111111111000000000000111111111111111111111111111111111111111111000000000001111100000000000011111111111111111111111111100000000000000000000000111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000001111111111111",
"1111110000000000000000000000000000000000000000000000001111111111111000000000000111111111111111111111111111111111111111111000000000001111100000000000001111111111111111111111111110000000000000000000001111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000011111111111111",
"1111110000000000000000000000000000000000000000000000011111111111111000000000000111111111111111111111111111111111111111110000000000011111110000000000001111111111111111111111111111000000000000000000001111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111100000000000000000000000000111111111111111",
"1111110000000000000000000000000000000000000000000001111111111111111000000000000111111111111111111111111111111111111111110000000000011111110000000000000111111111111111111111111111100000000000000000011111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000011111111111111111",
"1111110000000000000000000000000000000000000000001111111111111111111000000000000111111111111111111111111111111111111111100000000000111111111000000000000111111111111111111111111111100000000000000000111111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000111111111111111111",
"1111110000000000000000000000000000000000001111111111111111111111111000000000000111111111111111111111111111111111111111100000000000111111111000000000000011111111111111111111111111110000000000000001111111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000011111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111000000000001111111111100000000000011111111111111111111111111111000000000000001111111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111000000000001111111111100000000000001111111111111111111111111111000000000000011111111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111110000000000001111111111100000000000001111111111111111111111111111100000000000011111111111111111111111000000000000000000000000000000000111111111111111111100000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111000111111111111111111100000000000001111111110000000000000111111111111111111111111111111111111111111111000000000000000000000001111111111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111100000000000000000000000000000000000000111111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111100111111111111111111100000000000011111111111000000000000011111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111111111111111111111111100000000000011111111111000000000000001111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111000000000000000000000000000000000000000011111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111111111111111111111111100000000000011111111111100000000000001111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111111111111111111111111100000000000011111111111110000000000000111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111111111111111111111111100000000000011111111111110000000000000011111111111111111111111111111111111110000000000000000111111111111111111111111111111100011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111110011111110000000000000000000000000000000000000000000111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111111111111111001111111100000000000011111111111111000000000000011111111111111111111111111111111111100000000000000011111111111111111111111111111111000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111110001111100000000000001111111111111111110000000000000111111111111111111111111100000000000011111111111111111111111000000000000011111111111111111111111111111000111111100000000000011111111111111100000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000111111111111111111111111100001111100000000000011111111111111111111000000000000011111111111111111111111100000000000011111111111111111111111000000000000011111111111111111111111111110000111111100000000000011111111111111110000000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000001111100000000000111111111111111111111000000000000011111111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000000000000111111100000000000011111111111111110000000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000001111000000000000111111111111111111111100000000000001111111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000000000000111111100000000000011111111111111111000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000001111000000000001111111111111111111111100000000000001111111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000000000000111111100000000000011111111111111111100000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000001110000000000001111111111111111111111110000000000000111111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000000000000111111100000000000011111111111111111100000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000001100000000000011111111111111111111111110000000000000011111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000000000000111111100000000000011111111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1111110000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000001100000000000011111111111111111111111110000000000000011111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000000000000111111100000000000001111111111111111110000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1111100000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000001000000000000001111111111111111111111100000000000000000111111111111111111000000000000001111111111111111111110000000000000000000000000000000000000000000000111111000000000000001111111111111111110000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1110000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000001111111111111100000000000000000111111111111111111100000000000000000000000000000000000000000000000111110000000000000000011111111111111000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1110000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000001111111111111100000000000000000111111111111111111100000000000000000000000000000000000000000000000111110000000000000000011111111111111000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1111000000000000000001111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000011111111111111110000000000000000111111111111111111100000000000000000000000000000000000000000000000111110000000000000000011111111111111100000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111000011111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111100011111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111100000000000000000111111111111111111110000000000000000001111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111000000000000000011111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111000000000000000011111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111000000000000000001111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111100000000000000111111111111111111110000000000000000001111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111100000000000000111111111111111111110000000000000000001111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111110000000000000011111111111111111110000000000000000000111111111111111111000000000000001111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111110000000000000011111111111111111100000000000000000000111111111111111111000000000000011111111111111111111111000000000000000000001111111111111111111111000000000000000000111111111111111111100000000000000000111111111111111111111111111111110000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111000000000000001111111111111111100000000000000000000111111111111111110000000000000011111111111111111111000000000000000000000000011111111111111111111000000000000000000111111111111111111100000000000000000111111111111111111111111111111111000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111000000000000001111111111111111000000000000000000000011111111111111110000000000000111111111111111111100000000000000000000000000000111111111111111111000000000000000000111111111111111111110000000000000000111111111111111111111111111111111000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111000000000000001111111111111111000000000000000000000011111111111111110000000000000111111111111111111000000000000000000000000000000011111111111111111110000000000000001111111111111111111111100000000000011111111111111111111111111111111111000000000001111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111100000000000000111111111111111000000000000000000000001111111111111100000000000000111111111111111100000000000000000000000000000000000111111111111111110000000000000001111111111111111111111100000000000111111111111111111111111111111111111000000000001111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111100000000000000111111111111110000000000000000000000001111111111111100000000000001111111111111111000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111100000000000111111111111111111111111111111111111000000000001111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110000000000000111111111111110000000000000000000000001111111111111100000000000001111111111111110000000000000000000000000000000000000001111111111111110000000000000000011111111111111111111100000000000111111111111111111111111111111111111000000000001111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110000000000000011111111111110000000000000000000000000111111111111000000000000001111111111111100000000000000000000000000000000000000000011111111111110000000000000000001111111111111111111100000000000111111111111111111111111111111111111000000000011111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110000000000000011111111111100000000000000000000000000111111111111000000000000011111111111111000000000000000000000000000000000000000000001111111111110000000000000000000111111111111111111100000000000111111111111111111111111111111111111000000000011111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111000000000000011111111111100000000000010000000000000111111111111000000000000011111111111110000000000000000000111111110000000000000000001111111111110000000000000000000011111111111111111100000000000111111111111111111111111111111111111000000000011111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111000000000000001111111111000000000000011000000000000011111111110000000000000111111111111110000000000000000111111111111110000000000000000111111111110000000000000000000001111111111111111100000000000111111111111111111111111111111111111100000000011111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111100000000000001111111111000000000000111000000000000011111111110000000000000111111111111100000000000000011111111111111111100000000000000011111111110000000000000000000000111111111111111100000000000111111111111111111111111111111111111100000000011111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111100000000000001111111111000000000000111000000000000001111111100000000000000111111111111000000000000000111111111111111111110000000000000011111111110000000000000000000000011111111111111100000000000111111111111111111111111111111111111100000000011111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111100000000000000111111110000000000000111100000000000001111111100000000000001111111111111000000000000001111111111111111111111000000000000001111111110000000000000000000000001111111111111100000000000111111111111111111111111111111111111100000000011111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111110000000000000111111110000000000001111100000000000001111111100000000000001111111111111000000000000011111111111111111111111100000000000001111111110000000000000000000000000111111111111100000000000111111111111111111111111111111111111100000000011111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111110000000000000011111100000000000001111110000000000000111111000000000000011111111111110000000000000011111111111111111111111100000000000000111111110000000000000000000000000011111111111100000000000111111111111111111111111111111111111100000000011111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111110000000000000011111100000000000001111110000000000000111111000000000000011111111111110000000000000111111111111111111111111110000000000000111111110000000000000000000000000001111111111100000000000111111111111111111111111111111111111100000000111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111000000000000011111100000000000011111110000000000000111111000000000000011111111111110000000000000111111111111111111111111110000000000000111111110000000000000000000000000000111111111100000000000111111111111111111111111111111111111100000000111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111000000000000001111000000000000011111111000000000000011110000000000000111111111111110000000000001111111111111111111111111111000000000000111111110000000000001000000000000000011111111100000000000111111111111111111111111111111111111110000000111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111100000000000001111000000000000111111111000000000000011110000000000000111111111111100000000000001111111111111111111111111111000000000000011111110000000000001100000000000000001111111100000000000111111111111111111111111111111111111110000000111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111100000000000001111000000000000111111111000000000000011110000000000001111111111111100000000000001111111111111111111111111111000000000000011111110000000000001110000000000000000111111100000000000111111111111111111111111111111111111110000000111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111100000000000000110000000000000111111111100000000000001100000000000001111111111111100000000000001111111111111111111111111111000000000000011111110000000000001111000000000000000011111100000000000111111111111111111111111111111111111110000000111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111110000000000000110000000000001111111111100000000000001100000000000001111111111111100000000000001111111111111111111111111111000000000000011111110000000000001111100000000000000001111100000000000111111111111111111111111111111111111110000000111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111110000000000000100000000000001111111111110000000000000000000000000011111111111111100000000000001111111111111111111111111111000000000000011111110000000000001111110000000000000001111100000000000111111111111111111111111111111111111100000000111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111110000000000000000000000000011111111111111100000000000001111111111111111111111111111000000000000011111110000000000001111111000000000000000111100000000000111111111111111111111111111111111110000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000011111111111110000000000000000000000000011111111111111100000000000001111111111111111111111111111000000000000011111110000000000001111111100000000000000011100000000000111111111111111111111111111111111110000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111000000000000000000000000111111111111111110000000000001111111111111111111111111111000000000000011111110000000000001111111110000000000000001100000000000111111111111111111111111111111111110000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000111111111111111000000000000000000000000111111111111111110000000000001111111111111111111111111111000000000000111111110000000000001111111111000000000000000100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000111111111111111111111111110000000000000111111110000000000001111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000111111111111111111111111110000000000000111111110000000000001111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000011111111111111111111111100000000000000111111110000000000001111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111110000000000000000000011111111111111111111000000000000001111111111111111111111100000000000001111111110000000000001111111111111100000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111110000000000000000000011111111111111111111000000000000001111111111111111111111000000000000001111111110000000000001111111111111110000000000000000000000111111111111111111111111111111111111111100001111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111110000000000000000000111111111111111111111100000000000000111111111111111111110000000000000011111111110000000000001111111111111111000000000000000000000111111111111111111111111111111111111100000000011111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111000000000000000000111111111111111111111100000000000000001111111111111111000000000000000011111111110000000000001111111111111111100000000000000000000111111111111111111111111111111111111000000000001111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111000000000000000000111111111111111111111110000000000000000011111111111100000000000000000111111111110000000000001111111111111111110000000000000000000111111111111111111111111111111111110000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111000000000000000001111111111111111111111111000000000000000000011111100000000000000000000111111111110000000000001111111111111111111000000000000000000111111111111111111111111111111111110000000000000111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111100000000000000001111111111111111111111111100000000000000000000000000000000000000000001111111111110000000000001111111111111111111100000000000000000111111111111111111111111111111111100000000000000111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111100000000000000001111111111111111111111111110000000000000000000000000000000000000000011111111111110000000000001111111111111111111110000000000000000111111111111111111111111111111111100000000000000011111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111110000000000000011111111111111111111111111111000000000000000000000000000000000000000111111111111110000000000001111111111111111111111000000000000000111111111111111111111111111111111100000000000000011111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111110000000000000011111111111111111111111111111100000000000000000000000000000000000001111111111111110000000000001111111111111111111111100000000000000111111111111111111111111111111111100000000000000011111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111110000000000000011111111111111111111111111111110000000000000000000000000000000000011111111111111110000000000001111111111111111111111110000000000000111111111111111111111111111111111100000000000000111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111100000000000000001111111111111111111111111111111100000000000000000000000000000001111111111111111110000000000001111111111111111111111110000000000000011111111111111111111111111111111110000000000000111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111110000000000000000000011111111111111111111111111111111000000000000000000000000000111111111111111111000000000000000011111111111111111111000000000000000000111111111111111111111111111111110000000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111110000000000000000000011111111111111111111111111111111110000000000000000000000011111111111111111111000000000000000011111111111111111111000000000000000000111111111111111111111111111111111000000000001111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111110000000000000000000111111111111111111111111111111111111100000000000000000011111111111111111111111000000000000000011111111111111111111100000000000000000111111111111111111111111111111111100000000111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",			 
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");				

gameLabelVisible <= '1' when ((vPos >= (VD / 2) - 138) and (vPos < (VD / 2) - 74) and
                        (hPos >= (HD / 2) - 200) and (hPos < (HD / 2) + 200) and de = '1' and current_state = MENU and gameLabel(vPos - 102)(hPos - 120) = '0') else
						  '0';
						  
logoVisible <= '1' when ((vPos >= (VD / 2) + 45) and (vPos < (VD / 2) + 210) and
                   (hPos >= (HD / 2) - 100) and (hPos <(HD / 2) + 100) and
                    logo(vPos - ((VD / 2) + 45))(hPos - ((HD / 2) - 100)) 
                    = '0' and current_state = MENU) else
						  '0';	

StartGameLabelVisible <= '1' when ((vPos >= (VD / 2) - 48) and (vPos < (VD / 2) ) and
                        (hPos >= (HD / 2) - 200) and (hPos < (HD / 2) + 200) and de = '1' and current_state =  MENU  and StartGameLabel(vPos - 192)(hPos - 120) = '0' and label_delay_on = '1') else
						  '0';
p1_label_visible <= '1' when ((hPos > 100) and (hPos < 178) and (vPos > 446) and (vPos < 460) and de = '1' and p1_label(vPos-446)(hPos-100) = '0') else
							  '0';

p2_label_visible <= '1' when ((hPos > 450) and (hPos < 528) and (vPos > 446) and (vPos < 460) and de = '1' and p2_label(vPos-446)(hPos-450) = '0') else
							  '0';
	
						  
label_0p1_visible <= '1' when ((hPos > 141) and (hPos < 225) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_0(vPos-((VD/2)-62))(hPos-141) = '0' and (score_p1 = 0)) else
							  '0';						 
							 
label_1p1_visible <= '1' when ((hPos > 141) and (hPos < 225) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_1(vPos-((VD/2)-62))(hPos-141) = '0' and (score_p1 = 1)) else
							  '0';	
							 
label_2p1_visible <= '1' when ((hPos > 141) and (hPos < 225) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_2(vPos-((VD/2)-62))(hPos-141) = '0' and (score_p1 = 2)) else
							  '0';	

label_3p1_visible <= '1' when ((hPos > 141) and (hPos < 225) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_3(vPos-((VD/2)-62))(hPos-141) = '0' and (score_p1 = 3)) else
							  '0';

label_0p2_visible <= '1' when ((hPos > (HD-225)) and (hPos < (HD-141)) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_0(vPos-((VD/2)-62))(hPos-(HD-225)) = '0' and (score_p2 = 0)) else
							  '0';	
							  
label_1p2_visible <= '1' when ((hPos > (HD-225)) and (hPos < (HD-141)) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_1(vPos-((VD/2)-62))(hPos-(HD-225)) = '0' and (score_p2 = 1)) else
							  '0';	
							 
label_2p2_visible <= '1' when ((hPos > (HD-225)) and (hPos < (HD-141)) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_2(vPos-((VD/2)-62))(hPos-(HD-225)) = '0' and (score_p2 = 2)) else
							  '0';	

label_3p2_visible <= '1' when ((hPos > (HD-225)) and (hPos < (HD-141)) and (vPos > (VD/2)-62) and (vPos < (VD/2)+62) and de = '1' and label_3(vPos-((VD/2)-62))(hPos-(HD-225)) = '0' and (score_p2 = 3)) else
							  '0';

P1_Won_Label_visible <= '1' when ((hPos > 120) and (hPos < 520) and (vPos > 153) and (vPos < 327) and de = '1' and P1_Won_Label(vPos-153)(hPos-120) = '0' and current_state = P1_WIN) else
							  '0';		

P2_Won_Label_visible <= '1' when ((hPos > 120) and (hPos < 520) and (vPos > 153) and (vPos < 327) and de = '1' and P2_Won_Label(vPos-153)(hPos-120) = '0' and current_state = P2_WIN) else
							  '0';			  
							  

-- outputs
VGA_SYNC_N <= '0';
VGA_CLK <= clk25;

clk_div:process(CLOCK_50)
begin
    if(CLOCK_50'event and CLOCK_50 = '1')then
        clk25 <= not clk25;
    end if;
end process;

Horizontal_position_counter:process(clk25, RST)
begin
    if(RST = '0')then
        hpos <= 0;
    elsif(clk25'event and clk25 = '1')then
        if (hPos = (HD + HFP + HSP + HBP - 1)) then
            hPos <= 0;
        else
            hPos <= hPos + 1;
        end if;
    end if;
end process;

Vertical_position_counter:process(clk25, RST)
begin
    if(RST = '0')then
        vPos <= 0;
    elsif(clk25'event and clk25 = '1')then
        if(hPos = (HD + HFP + HSP + HBP - 1)) then
            if (vPos = (VD + VFP + VSP + VBP - 1)) then
                vPos <= 0;
            else
                vPos <= vPos + 1;
            end if;
        end if;
    end if;
end process;

Horizontal_Synchronisation:process(clk25, RST)
begin
    if(RST = '0')then
        hs    <= '0';
        VGA_HS <= '0';
    elsif(clk25'event and clk25 = '1')then
        if((hPos >= (HD + HFP)) AND (hPos < HD + HFP + HSP))then
            hs <= '0';
        else
            hs <= '1';
        end if;
        VGA_HS <= hs; -- delay one clock to account for pixel data delay
    end if;
end process;

Vertical_Synchronisation:process(clk25, RST)
begin
    if(RST = '0')then
        vs    <= '0';
        VGA_VS <= '0';
    elsif(clk25'event and clk25 = '1')then
        if((vPos >= (VD + VFP)) AND (vPos < VD + VFP + VSP))then
            vs <= '0';
        else
            vs <= '1';
        end if;
        VGA_VS <= vs; -- delay one clock to account for pixel data delay
    end if;
end process;

video_on:process(clk25, RST)
begin
    if(RST = '0')then
        de    <= '0';
        VGA_BLANK_N <= '0';
    elsif(clk25'event and clk25 = '1')then
        if(hPos < HD and vPos < VD)then
            de <= '1';
        else
            de <= '0';
        end if;
        VGA_BLANK_N <= de; -- delay one clock to align with pixel data
    end if;
end process;

draw:process(clk25, RST)
begin
	if(RST = '0')then
		VGA_R <= (others => '0');
      VGA_G <= (others => '0');
      VGA_B <= (others => '0');
	elsif(clk25'event and clk25 = '1')then
      if(de = '1')then
			if (current_state = MENU) then
				if (logoVisible = '1') then
					VGA_R <= "01011111";
					VGA_G <= (others => '0');
					VGA_B <= (others => '0');
				elsif (gameLabelVisible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif(StartGameLabelVisible = '1') then
					VGA_R <= (others => '1');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');					
				else
					VGA_R <= (others => '0');
					VGA_G <= (others => '0');
					VGA_B <= (others => '0');
				end if;
			elsif ((current_state = GAME) or (current_state = INITIAL)) then
				if ((hPos > p1_x1 and hPos < p1_x2) and (vPos > p1_y1 and vPos < p1_y2)) then
					VGA_R <= (others => '1');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif ((hPos > p2_x1 and hPos < p2_x2) and (vPos > p2_y1 and vPos < p2_y2)) then
					VGA_R <= (others => '1');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif ((hPos > ball_x1 and hPos < ball_x2) and (vPos > ball_y1 and vPos < ball_y2)) then
					VGA_R <= (others => '1');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_0p1_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_1p1_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_2p1_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_3p1_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_0p2_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_1p2_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_2p2_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif (label_3p2_visible = '1') then
					VGA_R <= (others => '0');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif(p1_label_visible = '1') then
					VGA_R <= (others => '1');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');
				elsif(p2_label_visible = '1') then
					VGA_R <= (others => '1');
					VGA_G <= (others => '1');
				   VGA_B <= (others => '1');					
				else
					VGA_R <= (others => '0');
					VGA_G <= (others => '0');
					VGA_B <= (others => '0');
				end if;  
			
			elsif((current_state = P1_WIN) or (current_state = P2_WIN)) then
				if (P1_Won_Label_visible = '1' or P2_Won_Label_visible = '1') then
					VGA_R <= (others => '1');
					VGA_G <= (others => '1');
					VGA_B <= (others => '1');	
				else
					VGA_R <= (others => '0');
					VGA_G <= (others => '0');
					VGA_B <= (others => '0');
				end if;
			end if;	
		else
			VGA_R <= (others => '0');
			VGA_G <= (others => '0');
			VGA_B <= (others => '0');
		end if;
   end if;
end process;

player1_move:process(clk25)
variable p1_move : std_logic_vector(0 to 1);
begin
	p1_move := p1_up & p1_down;
	if (clk25'event and clk25 = '1') then
		if (delayCounter1 = 50000) then
			delayCounter1 <= 0;
			case p1_move is
				when "10" =>
					if (p1_y2 < 480) then
						p1_y1 <= p1_y1 + 1;
						p1_y2 <= p1_y2 + 1;
					end if;
				when "01" =>
					if (p1_y1 > 0) then
						p1_y1 <= p1_y1 - 1;
						p1_y2 <= p1_y2 - 1;
					end if;
				when others =>
			end case;
		elsif(delayCounter2 = 50000 and current_state = INITIAL) then
			p1_x1 <= 20;
			p1_x2 <= 32;
			p1_y1 <= 195;
			p1_y2 <= 285;		
		else
			delayCounter1 <= delayCounter1 + 1;
		end if;
	end if;
end process;

player2_move:process(clk25)
variable p2_move : std_logic_vector(0 to 1);
begin
	p2_move := p2_up & p2_down;
	if (clk25'event and clk25 = '1') then
		if (delayCounter2 = 50000 and current_state = GAME) then
			delayCounter2 <= 0;
			case p2_move is
				when "10" =>
					if (p2_y2 < 480) then
						p2_y1 <= p2_y1 + 1;
						p2_y2 <= p2_y2 + 1;
					end if;		
				when "01" =>
					if (p2_y1 > 0) then
						p2_y1 <= p2_y1 - 1;
						p2_y2 <= p2_y2 - 1;
					end if;
				when others =>
			end case;
		elsif(delayCounter2 = 50000 and current_state = INITIAL) then
			p2_x1 <= 608;
			p2_x2 <= 620;
			p2_y1 <= 195;
			p2_y2 <= 285;	
		else
			delayCounter2 <= delayCounter2 + 1;
		end if;
	end if;
end process;

ball_move:process(clk25)
begin
	if (clk25'event and clk25 = '1') then
		if (delayCounter3 = 90000 and current_state = GAME) then
			delayCounter3 <= 0;
			goal_flag <= '0';
			if(ball_y1 = 0) then
				ball_move_v <= (-1)*ball_move_v;
				ball_y1 <= ball_y1 + 1;
				ball_y2 <= ball_y2 + 1;
			elsif(ball_y2 = 480) then
				ball_move_v <= (-1)*ball_move_v;
				ball_y2 <= ball_y2 - 1;
				ball_y1 <= ball_y1 - 1;
			elsif((ball_x2 = p2_x1) and (ball_y1 > p2_y1 and ball_y2 < p2_y2)) then
				ball_move_h <= (-1)*ball_move_h;
				ball_x2 <= ball_x2 - 1;
				ball_x1 <= ball_x1 - 1;
			elsif((ball_x1 = p1_x2) and (ball_y1 > p1_y1 and ball_y2 < p1_y2)) then
				ball_move_h <= (-1)*ball_move_h;
				ball_x2 <= ball_x2 + 1;
				ball_x1 <= ball_x1 + 1;
			elsif (ball_x2 = HD) then
				score_p1 <= score_p1 + 1;
				ball_x1 <= 313;
				ball_x2 <= 327;
				ball_y1 <= 233;
				ball_y2 <= 247;
				goal_flag <= '1';
			
				if(score_p1 = 3) then
					p1_w <= '1';
					p2_w <= '0';
				end if;
			elsif (ball_x1 = 0) then
				score_p2 <= score_p2 + 1;
				ball_x1 <= 313;
				ball_x2 <= 327;
				ball_y1 <= 233;
				ball_y2 <= 247;
				goal_flag <= '1';
				if(score_p2 = 3) then
					p1_w <= '0';
					p2_w <= '1';
				end if;
			else
				ball_y1 <= ball_y1 + ball_move_v;
				ball_y2 <= ball_y2 + ball_move_v;
				ball_x1 <= ball_x1 + ball_move_h;
				ball_x2 <= ball_x2 + ball_move_h;
			end if;	
		elsif(delayCounter3 = 90000 and current_state = INITIAL) then
			ball_x1 <= 313;
			ball_x2 <= 327;
			ball_y1 <= 233;
			ball_y2 <= 247;
		elsif(delayCounter3 = 90000 and (current_state = P1_WIN or current_state = P2_WIN)) then
			score_p1 <= 0;
			score_p2 <= 0;
			p1_w <= '0';
			p2_w <= '0';
		else
			delayCounter3 <= delayCounter3 + 1;
		end if;
	end if;
end process;


state_update : process(clk25,RST)
begin
	if (RST = '0') then
		current_state <= MENU;
	--	score_p1 <= 0;
	--	score_p2 <= 0;
	--	p1_w <= '0';
	--	p2_w <= '0';
	--	
	elsif (clk25'event and clk25 = '1') then
		current_state <= next_state;
	end if;
end process;

com_state : process(SW2, current_state)
begin
	case (current_state) is
		when (MENU) =>	
			if (SW2 = '1') then
				next_state <= MENU;
			else
				next_state <= INITIAL;
			end if;
		when (INITIAL) =>
			if((p1_up = '0' or p1_down = '0' or p2_up = '0' or p2_down = '0') and SW2 = '0') then
				next_state <= GAME;
			elsif(SW2 = '1') then
				next_state <= MENU;
			elsif(p1_w = '1') then
				next_state <= P1_WIN;
			elsif(p2_w = '1') then
				next_state <= P2_WIN;
			end if;
			
		when (GAME) =>
			if(goal_flag = '1') then
				next_state <= INITIAL;
				
			elsif (p1_w = '1' and p2_w = '0' and SW2 = '0') then
				next_state <= P1_WIN;
			elsif (p2_w = '1' and SW2 = '0' and p1_w = '0') then
				next_state <= P2_WIN;
			elsif (SW2 = '1') then
				next_state <= MENU;
			end if;
		when P1_WIN =>
			if(SW2 = '1') then
				next_state <= MENU;
			end if;
			
		when P2_WIN =>
			if(SW2 = '1') then
				next_state <= MENU;
			end if;
			
		end case;
end process;


delay : process(CLOCK_50)
begin
	if (CLOCK_50'event and CLOCK_50 = '1') then
		delay_label <= delay_label + 1;
		if(25_000_000 < delay_label and delay_label < 50_000_000) then
			label_delay_on <= '1';
		elsif(delay_label < 25_000_000) then
			label_delay_on <= '0';
		elsif(delay_label = 50_000_000) then
			delay_label <= 0;
		end if;
	end if;
end process;





end;